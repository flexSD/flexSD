library verilog;
use verilog.vl_types.all;
entity UDFDL5E_UDP_X is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end UDFDL5E_UDP_X;
