library verilog;
use verilog.vl_types.all;
entity sinegen_tb is
end sinegen_tb;
