library verilog;
use verilog.vl_types.all;
entity lut_mux4 is
    // This module cannot be connected to from
    // VHDL because it has unnamed ports.
end lut_mux4;
