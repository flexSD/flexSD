`timescale 100ps/1ps

/* 24 bit second order 10x virtualized Sigma Delta modulator 
 * 
 * flexSD project
 * Dan Kouba, 2012
 * 
 * CURRENT LIMITATIONS (6/7/12) :
 * Sigma delta assumes that slice is only implementing one filter of arbitrary order, with hardware inputs and outputs (aka no other filters before or after)
 *    - Cannot log multiple values within one slice run
 *    - 
 */
 
module second_order_sigdel_virtualized(
  
  clock_200,
  clock_20,
  reset,
  mod_enable,
  
  write_address_in,
  write_enable_in,
  
  log_address,
  log_value_reconstructed,  
  log_bitstream,
  
  input_data,
  virtualized_bitstream_reg,
  
  external_bitstreams_in,
  external_bitstream_address,
  external_bitstream_reg

  
);

/* Internal prameters */
parameter input_bitwidth          = 24;
parameter accumulator_bitwidth    = 36;

/* Define full scale positive and negative values for the feedback loop
 * These values are full scale values as wide as the input bitwidth, sign extended to the accumulator's bitwidth */
`define full_neg {{(accumulator_bitwidth - input_bitwidth + 1){1'b1}}, {(input_bitwidth-1){1'b0}}}
`define full_pos {{(accumulator_bitwidth - input_bitwidth + 1){1'b0}}, {(input_bitwidth-1){1'b1}}}

/* Module inputs and outputs */
input                      clock_200, clock_20;
input                      reset;
input                      mod_enable;                                    // Enables whole modulator

input          [3:0]       write_address_in;                              // Address for input value storage RAM
input                      write_enable_in;                               // Enable for writing new value to input value storage RAM

input          [3:0]       log_address;                                   // Address of the bitstream to log (0-9)
output         [23:0]      log_value_reconstructed;                       // Reconstructed value of the logged bitstream
output                     log_bitstream;                                 // Bitstream that has been logged, USED AS FEEDBACK SIGMA DELTA STREAM FOR SLICE!!!!!

input   signed [23:0]      input_data;                                    // Input to the value storage ram front end
output         [9:0]       virtualized_bitstream_reg;                     // 10 bit register containing all bitstreams from the virtual modulators

input          [3:0]       external_bitstreams_in;                        // Input bitstreams from ADC - synchronized with the output bitstream register
input          [1:0]       external_bitstream_address;                    // Address of external bitstream to output to the storage register
output                     external_bitstream_reg;                        // Register that contains external ADCs bitstreams, synced with virtualized bitstream register

/* Internal wires and registers */
wire    signed [accumulator_bitwidth - 1:0]      fb;                      // Feedback signal, 28 bits, but only holds a 24 bit full scale number as defined by the parameters above
wire    signed [accumulator_bitwidth - 1:0]      error_1;                 // First error signal, equals input minus the feedback signal
wire    signed [accumulator_bitwidth - 1:0]      error_2;                 // Second error signal, equals the output of the nondelaying integrator minus the feedback signal
wire    signed [accumulator_bitwidth - 1:0]      adder_1_out;             // Adder that creates the nondelaying integrator
wire    signed [accumulator_bitwidth - 1:0]      accumulator_1_out;       // Nondelaying integrator's z^-1 block
wire    signed [accumulator_bitwidth - 1:0]      accumulator_2_out;       // Delaying integrator's z^-1 block
wire                                             comp_out;                // Output of the comparator, also the output bitstream

// For RAM addressing
reg            [1:0]                             mod_enable_delay_reg;    // Write addresses are one clock behind the read addresses (due to reg on output of accumulator RAM)
reg            [3:0]                             address_counter;         // Address counter for read and write addresses
reg            [3:0]                             address_delay_reg;       // Delay the address counter value one clock from the read cycle for the write cycle
wire    signed [23:0]                            value_storage_out;       // Output of the value storage RAM
reg                                              log_bitstream_i;         // Addressed bit of the output bitstream register to log and reconstruct
//reg            [3:0]                             log_address_reg;         // Clocks in new address to log when the logging trigger comes in
wire           [3:0]                             acc_read_adr;            // Accumulator read address, generated by internal counter
wire           [3:0]                             acc_write_adr;           // Accumulator write address, generated from delayed read address

/* Address Counter */

// Instantiate counter - counts from 0 to 9 and then loops
always@(negedge clock_200) begin
  
  if(reset) address_counter = 4'd9;       // Always start at address '0' after reset
  else if(mod_enable) begin
    
    if(address_counter == 4'd9) address_counter <= 4'b0;    // Reset to 0 if at maximum count (9)
    else address_counter <= address_counter + 1'b1;         // Otherwise add 1 to current count
    
  end
  
end

/* Enable Delay Alignment */

always@(negedge clock_200) begin
  
  if(reset) begin
  
    mod_enable_delay_reg <= 2'b0;
    address_delay_reg <= 4'b0;
  
  end else begin  
    
    // Create delayed enable signal for write back operations
    mod_enable_delay_reg[1] <= mod_enable_delay_reg[0];
    mod_enable_delay_reg[0] <= mod_enable;  
    
    // Create delayed address for write back operation (delayed one clock)
    address_delay_reg <= address_counter;
    
  end
  
end

// Address assigns
assign acc_read_adr = address_counter;
assign acc_write_adr = address_delay_reg;

// Enable assigns
assign acc_read_en = mod_enable_delay_reg[0];
assign acc_write_en = mod_enable_delay_reg[1];

lattice_ram_24bit_16word value_storage_ram(

  .WrAddress(write_address_in), 
  .Data(input_data), 
  .WrClock(clock_200), 
  .WE(write_enable_in), 
  .WrClockEn(write_enable_in), 
  .RdAddress(acc_read_adr),
  .RdClock(clock_200),
  .RdClockEn(acc_read_en),
  .Reset(reset),
  .Q(value_storage_out)

);

lattice_ram_36bit_16 accumulator_1(

  .WrAddress(acc_write_adr), 
  .Data(adder_1_out), 
  .WrClock(clock_200), 
  .WE(acc_write_en), 
  .WrClockEn(acc_write_en), 
  .RdAddress(acc_read_adr),
  .RdClock(clock_200),
  .RdClockEn(acc_read_en),
  .Reset(reset),
  .Q(accumulator_1_out)

);

lattice_ram_36bit_16 accumulator_2(

  .WrAddress(acc_write_adr), 
  .Data(accumulator_2_out + error_2), 
  .WrClock(clock_200), 
  .WE(acc_write_en), 
  .WrClockEn(acc_write_en), 
  .RdAddress(acc_read_adr),
  .RdClock(clock_200),
  .RdClockEn(acc_read_en),
  .Reset(reset),
  .Q(accumulator_2_out)

);

reconstruction_filter recon_filter(
  .clock(clock_20),
  .reset(reset),
  .bitstream_in(log_bitstream),
  .out(log_value_reconstructed)
  
);

/* Bitstream Storage */

// Create shift register on output that shifts in each bit as it is created by the virtualized modulators
reg     [9:0]      bitstream_reg_i;                 // Internal bitstream register
reg     [9:0]      virtualized_bitstream_reg_i;     // Register retains the last 10 sigma delta output bits for the slice to use in its virtual cycles
reg     [3:0]      external_bitstream_in_i;         // Stores external bitstream values from ADC at same interval as the virtualized bitstream register
reg                external_bitstream_reg_i;        // Stores external bitstream value chosen by external bitstream address

always@(posedge clock_200) begin
  
  if(reset) begin
  
    bitstream_reg_i <= 10'b0;
    virtualized_bitstream_reg_i <= 10'b0;
    external_bitstream_in_i <= 4'b0;
    external_bitstream_reg_i <= 1'b0;
  
  end else if(mod_enable_delay_reg[0]) begin    // Must be delayed one from the modulator enable so that the ram can read out and adds can happen before the bitstream is written
  
    bitstream_reg_i <= { comp_out, bitstream_reg_i[9:1] };
    
    /* Every 10th cycle copy shift register data to external register - outputted to slice
     *sim:/slice_vliw_sigdel_tb/slice1/add_sub_result_B

     * mod_enable_delay_reg[1] check is there to prevent clock in of bitstream data on initialization of the modulator.
     * This prevents uninitialized data from being clocked into the filter when it is started up and ensures a register full of zeros at the beginning.
     * 
     * Addressing:
     * [9:0]   - Internal virtual sigma delta bitstreams, addressed in order of slice operation (address 0 is the first order of the slice)
     * [13:10] - External ADC bitstreams, synchronized to this clock domain
     */
    if( (address_counter == 4'd0) && (mod_enable_delay_reg[1]) ) begin
       
       virtualized_bitstream_reg_i <= { comp_out, bitstream_reg_i[9:1] };      
       external_bitstream_in_i <= external_bitstreams_in[3:0];
       
    end
  
  end
  
end

assign virtualized_bitstream_reg = virtualized_bitstream_reg_i;

/* Logging handler */
/*
//limited to handling only one log per filter cycle!!!!!!!!!!  Multple logs will cause output of reconstruction filter to become nonsensical, as multiple signals would mix
always@(posedge clock_200) begin
  
  if(log_trigger) log_address_reg <= log_address;

end
 */   
// Continuously assinged mux: logging address is the select, bitstream reg bits are the inputs, logged bitstream is the output
always@(log_address or virtualized_bitstream_reg_i) begin

  case(log_address)
      
    default: log_bitstream_i <= virtualized_bitstream_reg_i[0];   // We only have 10 addresses to access, and 16 possible addresses so any invalid address results in the first bitstream
    4'd0:    log_bitstream_i <= virtualized_bitstream_reg_i[0];
    4'd1:    log_bitstream_i <= virtualized_bitstream_reg_i[1];
    4'd2:    log_bitstream_i <= virtualized_bitstream_reg_i[2];
    4'd3:    log_bitstream_i <= virtualized_bitstream_reg_i[3];
    4'd4:    log_bitstream_i <= virtualized_bitstream_reg_i[4];
    4'd5:    log_bitstream_i <= virtualized_bitstream_reg_i[5];
    4'd6:    log_bitstream_i <= virtualized_bitstream_reg_i[6];
    4'd7:    log_bitstream_i <= virtualized_bitstream_reg_i[7];
    4'd8:    log_bitstream_i <= virtualized_bitstream_reg_i[8];
    4'd9:    log_bitstream_i <= virtualized_bitstream_reg_i[9];
      
  endcase
    
end

assign log_bitstream = log_bitstream_i;

// Mux external bitstreams out to the external bitstream output based on address from VLIW
always@(external_bitstream_address or external_bitstream_in_i) begin
  
  case(external_bitstream_address)
    
    default:  external_bitstream_reg_i <= external_bitstream_in_i[0];
    2'd0:     external_bitstream_reg_i <= external_bitstream_in_i[0];
    2'd1:     external_bitstream_reg_i <= external_bitstream_in_i[1];
    2'd2:     external_bitstream_reg_i <= external_bitstream_in_i[2];
    2'd3:     external_bitstream_reg_i <= external_bitstream_in_i[3];
    
  endcase
  
end

assign external_bitstream_reg = external_bitstream_reg_i;

/* Adders, output comparator and signal routing */

assign adder_1_out = accumulator_1_out + error_1;
assign comp_out = !accumulator_2_out[accumulator_bitwidth - 1];  // To do comparison, grab sign bit and invert (due to 2's complement)

assign error_1 = value_storage_out - fb;
assign error_2 = adder_1_out - fb;

assign fb = comp_out ? `full_pos : `full_neg;          //Comparator, 24 bit full scale output

endmodule