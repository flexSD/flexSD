library verilog;
use verilog.vl_types.all;
entity OB is
    port(
        I               : in     vl_logic;
        O               : out    vl_logic
    );
end OB;
