library verilog;
use verilog.vl_types.all;
entity state_ram_tb is
end state_ram_tb;
