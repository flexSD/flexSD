library verilog;
use verilog.vl_types.all;
entity XOR11 is
    port(
        A               : in     vl_logic;
        B               : in     vl_logic;
        C               : in     vl_logic;
        D               : in     vl_logic;
        E               : in     vl_logic;
        F               : in     vl_logic;
        G               : in     vl_logic;
        H               : in     vl_logic;
        I               : in     vl_logic;
        J               : in     vl_logic;
        K               : in     vl_logic;
        Z               : out    vl_logic
    );
end XOR11;
