library verilog;
use verilog.vl_types.all;
entity sigdel_tb is
    generic(
        input_bitwidth  : integer := 12
    );
end sigdel_tb;
