library verilog;
use verilog.vl_types.all;
entity VLIW_tb is
end VLIW_tb;
