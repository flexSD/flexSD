library verilog;
use verilog.vl_types.all;
entity XOR21 is
    port(
        A               : in     vl_logic;
        B               : in     vl_logic;
        C               : in     vl_logic;
        D               : in     vl_logic;
        E               : in     vl_logic;
        F               : in     vl_logic;
        G               : in     vl_logic;
        H               : in     vl_logic;
        I               : in     vl_logic;
        J               : in     vl_logic;
        K               : in     vl_logic;
        L               : in     vl_logic;
        M               : in     vl_logic;
        N               : in     vl_logic;
        O               : in     vl_logic;
        P               : in     vl_logic;
        Q               : in     vl_logic;
        R               : in     vl_logic;
        S               : in     vl_logic;
        T               : in     vl_logic;
        U               : in     vl_logic;
        Z               : out    vl_logic
    );
end XOR21;
