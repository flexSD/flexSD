library verilog;
use verilog.vl_types.all;
entity GSR is
    port(
        GSR             : in     vl_logic
    );
end GSR;
