library verilog;
use verilog.vl_types.all;
entity MULT18X18ADDSUBSUMB is
    generic(
        REG_INPUTA0_CLK : string  := "NONE";
        REG_INPUTA0_CE  : string  := "CE0";
        REG_INPUTA0_RST : string  := "RST0";
        REG_INPUTA1_CLK : string  := "NONE";
        REG_INPUTA1_CE  : string  := "CE0";
        REG_INPUTA1_RST : string  := "RST0";
        REG_INPUTA2_CLK : string  := "NONE";
        REG_INPUTA2_CE  : string  := "CE0";
        REG_INPUTA2_RST : string  := "RST0";
        REG_INPUTA3_CLK : string  := "NONE";
        REG_INPUTA3_CE  : string  := "CE0";
        REG_INPUTA3_RST : string  := "RST0";
        REG_INPUTB0_CLK : string  := "NONE";
        REG_INPUTB0_CE  : string  := "CE0";
        REG_INPUTB0_RST : string  := "RST0";
        REG_INPUTB1_CLK : string  := "NONE";
        REG_INPUTB1_CE  : string  := "CE0";
        REG_INPUTB1_RST : string  := "RST0";
        REG_INPUTB2_CLK : string  := "NONE";
        REG_INPUTB2_CE  : string  := "CE0";
        REG_INPUTB2_RST : string  := "RST0";
        REG_INPUTB3_CLK : string  := "NONE";
        REG_INPUTB3_CE  : string  := "CE0";
        REG_INPUTB3_RST : string  := "RST0";
        REG_PIPELINE0_CLK: string  := "NONE";
        REG_PIPELINE0_CE: string  := "CE0";
        REG_PIPELINE0_RST: string  := "RST0";
        REG_PIPELINE1_CLK: string  := "NONE";
        REG_PIPELINE1_CE: string  := "CE0";
        REG_PIPELINE1_RST: string  := "RST0";
        REG_PIPELINE2_CLK: string  := "NONE";
        REG_PIPELINE2_CE: string  := "CE0";
        REG_PIPELINE2_RST: string  := "RST0";
        REG_PIPELINE3_CLK: string  := "NONE";
        REG_PIPELINE3_CE: string  := "CE0";
        REG_PIPELINE3_RST: string  := "RST0";
        REG_OUTPUT_CLK  : string  := "NONE";
        REG_OUTPUT_CE   : string  := "CE0";
        REG_OUTPUT_RST  : string  := "RST0";
        REG_SIGNEDA_0_CLK: string  := "NONE";
        REG_SIGNEDA_0_CE: string  := "CE0";
        REG_SIGNEDA_0_RST: string  := "RST0";
        REG_SIGNEDA_1_CLK: string  := "NONE";
        REG_SIGNEDA_1_CE: string  := "CE0";
        REG_SIGNEDA_1_RST: string  := "RST0";
        REG_SIGNEDB_0_CLK: string  := "NONE";
        REG_SIGNEDB_0_CE: string  := "CE0";
        REG_SIGNEDB_0_RST: string  := "RST0";
        REG_SIGNEDB_1_CLK: string  := "NONE";
        REG_SIGNEDB_1_CE: string  := "CE0";
        REG_SIGNEDB_1_RST: string  := "RST0";
        REG_ADDNSUB1_0_CLK: string  := "NONE";
        REG_ADDNSUB1_0_CE: string  := "CE0";
        REG_ADDNSUB1_0_RST: string  := "RST0";
        REG_ADDNSUB1_1_CLK: string  := "NONE";
        REG_ADDNSUB1_1_CE: string  := "CE0";
        REG_ADDNSUB1_1_RST: string  := "RST0";
        REG_ADDNSUB3_0_CLK: string  := "NONE";
        REG_ADDNSUB3_0_CE: string  := "CE0";
        REG_ADDNSUB3_0_RST: string  := "RST0";
        REG_ADDNSUB3_1_CLK: string  := "NONE";
        REG_ADDNSUB3_1_CE: string  := "CE0";
        REG_ADDNSUB3_1_RST: string  := "RST0";
        GSR             : string  := "ENABLED"
    );
    port(
        SUM37           : out    vl_logic;
        SUM36           : out    vl_logic;
        SUM35           : out    vl_logic;
        SUM34           : out    vl_logic;
        SUM33           : out    vl_logic;
        SUM32           : out    vl_logic;
        SUM31           : out    vl_logic;
        SUM30           : out    vl_logic;
        SUM29           : out    vl_logic;
        SUM28           : out    vl_logic;
        SUM27           : out    vl_logic;
        SUM26           : out    vl_logic;
        SUM25           : out    vl_logic;
        SUM24           : out    vl_logic;
        SUM23           : out    vl_logic;
        SUM22           : out    vl_logic;
        SUM21           : out    vl_logic;
        SUM20           : out    vl_logic;
        SUM19           : out    vl_logic;
        SUM18           : out    vl_logic;
        SUM17           : out    vl_logic;
        SUM16           : out    vl_logic;
        SUM15           : out    vl_logic;
        SUM14           : out    vl_logic;
        SUM13           : out    vl_logic;
        SUM12           : out    vl_logic;
        SUM11           : out    vl_logic;
        SUM10           : out    vl_logic;
        SUM9            : out    vl_logic;
        SUM8            : out    vl_logic;
        SUM7            : out    vl_logic;
        SUM6            : out    vl_logic;
        SUM5            : out    vl_logic;
        SUM4            : out    vl_logic;
        SUM3            : out    vl_logic;
        SUM2            : out    vl_logic;
        SUM1            : out    vl_logic;
        SUM0            : out    vl_logic;
        SROA17          : out    vl_logic;
        SROA16          : out    vl_logic;
        SROA15          : out    vl_logic;
        SROA14          : out    vl_logic;
        SROA13          : out    vl_logic;
        SROA12          : out    vl_logic;
        SROA11          : out    vl_logic;
        SROA10          : out    vl_logic;
        SROA9           : out    vl_logic;
        SROA8           : out    vl_logic;
        SROA7           : out    vl_logic;
        SROA6           : out    vl_logic;
        SROA5           : out    vl_logic;
        SROA4           : out    vl_logic;
        SROA3           : out    vl_logic;
        SROA2           : out    vl_logic;
        SROA1           : out    vl_logic;
        SROA0           : out    vl_logic;
        SROB17          : out    vl_logic;
        SROB16          : out    vl_logic;
        SROB15          : out    vl_logic;
        SROB14          : out    vl_logic;
        SROB13          : out    vl_logic;
        SROB12          : out    vl_logic;
        SROB11          : out    vl_logic;
        SROB10          : out    vl_logic;
        SROB9           : out    vl_logic;
        SROB8           : out    vl_logic;
        SROB7           : out    vl_logic;
        SROB6           : out    vl_logic;
        SROB5           : out    vl_logic;
        SROB4           : out    vl_logic;
        SROB3           : out    vl_logic;
        SROB2           : out    vl_logic;
        SROB1           : out    vl_logic;
        SROB0           : out    vl_logic;
        A017            : in     vl_logic;
        A016            : in     vl_logic;
        A015            : in     vl_logic;
        A014            : in     vl_logic;
        A013            : in     vl_logic;
        A012            : in     vl_logic;
        A011            : in     vl_logic;
        A010            : in     vl_logic;
        A09             : in     vl_logic;
        A08             : in     vl_logic;
        A07             : in     vl_logic;
        A06             : in     vl_logic;
        A05             : in     vl_logic;
        A04             : in     vl_logic;
        A03             : in     vl_logic;
        A02             : in     vl_logic;
        A01             : in     vl_logic;
        A00             : in     vl_logic;
        A117            : in     vl_logic;
        A116            : in     vl_logic;
        A115            : in     vl_logic;
        A114            : in     vl_logic;
        A113            : in     vl_logic;
        A112            : in     vl_logic;
        A111            : in     vl_logic;
        A110            : in     vl_logic;
        A19             : in     vl_logic;
        A18             : in     vl_logic;
        A17             : in     vl_logic;
        A16             : in     vl_logic;
        A15             : in     vl_logic;
        A14             : in     vl_logic;
        A13             : in     vl_logic;
        A12             : in     vl_logic;
        A11             : in     vl_logic;
        A10             : in     vl_logic;
        A217            : in     vl_logic;
        A216            : in     vl_logic;
        A215            : in     vl_logic;
        A214            : in     vl_logic;
        A213            : in     vl_logic;
        A212            : in     vl_logic;
        A211            : in     vl_logic;
        A210            : in     vl_logic;
        A29             : in     vl_logic;
        A28             : in     vl_logic;
        A27             : in     vl_logic;
        A26             : in     vl_logic;
        A25             : in     vl_logic;
        A24             : in     vl_logic;
        A23             : in     vl_logic;
        A22             : in     vl_logic;
        A21             : in     vl_logic;
        A20             : in     vl_logic;
        A317            : in     vl_logic;
        A316            : in     vl_logic;
        A315            : in     vl_logic;
        A314            : in     vl_logic;
        A313            : in     vl_logic;
        A312            : in     vl_logic;
        A311            : in     vl_logic;
        A310            : in     vl_logic;
        A39             : in     vl_logic;
        A38             : in     vl_logic;
        A37             : in     vl_logic;
        A36             : in     vl_logic;
        A35             : in     vl_logic;
        A34             : in     vl_logic;
        A33             : in     vl_logic;
        A32             : in     vl_logic;
        A31             : in     vl_logic;
        A30             : in     vl_logic;
        B017            : in     vl_logic;
        B016            : in     vl_logic;
        B015            : in     vl_logic;
        B014            : in     vl_logic;
        B013            : in     vl_logic;
        B012            : in     vl_logic;
        B011            : in     vl_logic;
        B010            : in     vl_logic;
        B09             : in     vl_logic;
        B08             : in     vl_logic;
        B07             : in     vl_logic;
        B06             : in     vl_logic;
        B05             : in     vl_logic;
        B04             : in     vl_logic;
        B03             : in     vl_logic;
        B02             : in     vl_logic;
        B01             : in     vl_logic;
        B00             : in     vl_logic;
        B117            : in     vl_logic;
        B116            : in     vl_logic;
        B115            : in     vl_logic;
        B114            : in     vl_logic;
        B113            : in     vl_logic;
        B112            : in     vl_logic;
        B111            : in     vl_logic;
        B110            : in     vl_logic;
        B19             : in     vl_logic;
        B18             : in     vl_logic;
        B17             : in     vl_logic;
        B16             : in     vl_logic;
        B15             : in     vl_logic;
        B14             : in     vl_logic;
        B13             : in     vl_logic;
        B12             : in     vl_logic;
        B11             : in     vl_logic;
        B10             : in     vl_logic;
        B217            : in     vl_logic;
        B216            : in     vl_logic;
        B215            : in     vl_logic;
        B214            : in     vl_logic;
        B213            : in     vl_logic;
        B212            : in     vl_logic;
        B211            : in     vl_logic;
        B210            : in     vl_logic;
        B29             : in     vl_logic;
        B28             : in     vl_logic;
        B27             : in     vl_logic;
        B26             : in     vl_logic;
        B25             : in     vl_logic;
        B24             : in     vl_logic;
        B23             : in     vl_logic;
        B22             : in     vl_logic;
        B21             : in     vl_logic;
        B20             : in     vl_logic;
        B317            : in     vl_logic;
        B316            : in     vl_logic;
        B315            : in     vl_logic;
        B314            : in     vl_logic;
        B313            : in     vl_logic;
        B312            : in     vl_logic;
        B311            : in     vl_logic;
        B310            : in     vl_logic;
        B39             : in     vl_logic;
        B38             : in     vl_logic;
        B37             : in     vl_logic;
        B36             : in     vl_logic;
        B35             : in     vl_logic;
        B34             : in     vl_logic;
        B33             : in     vl_logic;
        B32             : in     vl_logic;
        B31             : in     vl_logic;
        B30             : in     vl_logic;
        SRIA17          : in     vl_logic;
        SRIA16          : in     vl_logic;
        SRIA15          : in     vl_logic;
        SRIA14          : in     vl_logic;
        SRIA13          : in     vl_logic;
        SRIA12          : in     vl_logic;
        SRIA11          : in     vl_logic;
        SRIA10          : in     vl_logic;
        SRIA9           : in     vl_logic;
        SRIA8           : in     vl_logic;
        SRIA7           : in     vl_logic;
        SRIA6           : in     vl_logic;
        SRIA5           : in     vl_logic;
        SRIA4           : in     vl_logic;
        SRIA3           : in     vl_logic;
        SRIA2           : in     vl_logic;
        SRIA1           : in     vl_logic;
        SRIA0           : in     vl_logic;
        SRIB17          : in     vl_logic;
        SRIB16          : in     vl_logic;
        SRIB15          : in     vl_logic;
        SRIB14          : in     vl_logic;
        SRIB13          : in     vl_logic;
        SRIB12          : in     vl_logic;
        SRIB11          : in     vl_logic;
        SRIB10          : in     vl_logic;
        SRIB9           : in     vl_logic;
        SRIB8           : in     vl_logic;
        SRIB7           : in     vl_logic;
        SRIB6           : in     vl_logic;
        SRIB5           : in     vl_logic;
        SRIB4           : in     vl_logic;
        SRIB3           : in     vl_logic;
        SRIB2           : in     vl_logic;
        SRIB1           : in     vl_logic;
        SRIB0           : in     vl_logic;
        SIGNEDA         : in     vl_logic;
        SIGNEDB         : in     vl_logic;
        ADDNSUB1        : in     vl_logic;
        ADDNSUB3        : in     vl_logic;
        CE0             : in     vl_logic;
        CE1             : in     vl_logic;
        CE2             : in     vl_logic;
        CE3             : in     vl_logic;
        CLK0            : in     vl_logic;
        CLK1            : in     vl_logic;
        CLK2            : in     vl_logic;
        CLK3            : in     vl_logic;
        RST0            : in     vl_logic;
        RST1            : in     vl_logic;
        RST2            : in     vl_logic;
        RST3            : in     vl_logic;
        SOURCEA0        : in     vl_logic;
        SOURCEA1        : in     vl_logic;
        SOURCEA2        : in     vl_logic;
        SOURCEA3        : in     vl_logic;
        SOURCEB0        : in     vl_logic;
        SOURCEB1        : in     vl_logic;
        SOURCEB2        : in     vl_logic;
        SOURCEB3        : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of REG_INPUTA0_CLK : constant is 1;
    attribute mti_svvh_generic_type of REG_INPUTA0_CE : constant is 1;
    attribute mti_svvh_generic_type of REG_INPUTA0_RST : constant is 1;
    attribute mti_svvh_generic_type of REG_INPUTA1_CLK : constant is 1;
    attribute mti_svvh_generic_type of REG_INPUTA1_CE : constant is 1;
    attribute mti_svvh_generic_type of REG_INPUTA1_RST : constant is 1;
    attribute mti_svvh_generic_type of REG_INPUTA2_CLK : constant is 1;
    attribute mti_svvh_generic_type of REG_INPUTA2_CE : constant is 1;
    attribute mti_svvh_generic_type of REG_INPUTA2_RST : constant is 1;
    attribute mti_svvh_generic_type of REG_INPUTA3_CLK : constant is 1;
    attribute mti_svvh_generic_type of REG_INPUTA3_CE : constant is 1;
    attribute mti_svvh_generic_type of REG_INPUTA3_RST : constant is 1;
    attribute mti_svvh_generic_type of REG_INPUTB0_CLK : constant is 1;
    attribute mti_svvh_generic_type of REG_INPUTB0_CE : constant is 1;
    attribute mti_svvh_generic_type of REG_INPUTB0_RST : constant is 1;
    attribute mti_svvh_generic_type of REG_INPUTB1_CLK : constant is 1;
    attribute mti_svvh_generic_type of REG_INPUTB1_CE : constant is 1;
    attribute mti_svvh_generic_type of REG_INPUTB1_RST : constant is 1;
    attribute mti_svvh_generic_type of REG_INPUTB2_CLK : constant is 1;
    attribute mti_svvh_generic_type of REG_INPUTB2_CE : constant is 1;
    attribute mti_svvh_generic_type of REG_INPUTB2_RST : constant is 1;
    attribute mti_svvh_generic_type of REG_INPUTB3_CLK : constant is 1;
    attribute mti_svvh_generic_type of REG_INPUTB3_CE : constant is 1;
    attribute mti_svvh_generic_type of REG_INPUTB3_RST : constant is 1;
    attribute mti_svvh_generic_type of REG_PIPELINE0_CLK : constant is 1;
    attribute mti_svvh_generic_type of REG_PIPELINE0_CE : constant is 1;
    attribute mti_svvh_generic_type of REG_PIPELINE0_RST : constant is 1;
    attribute mti_svvh_generic_type of REG_PIPELINE1_CLK : constant is 1;
    attribute mti_svvh_generic_type of REG_PIPELINE1_CE : constant is 1;
    attribute mti_svvh_generic_type of REG_PIPELINE1_RST : constant is 1;
    attribute mti_svvh_generic_type of REG_PIPELINE2_CLK : constant is 1;
    attribute mti_svvh_generic_type of REG_PIPELINE2_CE : constant is 1;
    attribute mti_svvh_generic_type of REG_PIPELINE2_RST : constant is 1;
    attribute mti_svvh_generic_type of REG_PIPELINE3_CLK : constant is 1;
    attribute mti_svvh_generic_type of REG_PIPELINE3_CE : constant is 1;
    attribute mti_svvh_generic_type of REG_PIPELINE3_RST : constant is 1;
    attribute mti_svvh_generic_type of REG_OUTPUT_CLK : constant is 1;
    attribute mti_svvh_generic_type of REG_OUTPUT_CE : constant is 1;
    attribute mti_svvh_generic_type of REG_OUTPUT_RST : constant is 1;
    attribute mti_svvh_generic_type of REG_SIGNEDA_0_CLK : constant is 1;
    attribute mti_svvh_generic_type of REG_SIGNEDA_0_CE : constant is 1;
    attribute mti_svvh_generic_type of REG_SIGNEDA_0_RST : constant is 1;
    attribute mti_svvh_generic_type of REG_SIGNEDA_1_CLK : constant is 1;
    attribute mti_svvh_generic_type of REG_SIGNEDA_1_CE : constant is 1;
    attribute mti_svvh_generic_type of REG_SIGNEDA_1_RST : constant is 1;
    attribute mti_svvh_generic_type of REG_SIGNEDB_0_CLK : constant is 1;
    attribute mti_svvh_generic_type of REG_SIGNEDB_0_CE : constant is 1;
    attribute mti_svvh_generic_type of REG_SIGNEDB_0_RST : constant is 1;
    attribute mti_svvh_generic_type of REG_SIGNEDB_1_CLK : constant is 1;
    attribute mti_svvh_generic_type of REG_SIGNEDB_1_CE : constant is 1;
    attribute mti_svvh_generic_type of REG_SIGNEDB_1_RST : constant is 1;
    attribute mti_svvh_generic_type of REG_ADDNSUB1_0_CLK : constant is 1;
    attribute mti_svvh_generic_type of REG_ADDNSUB1_0_CE : constant is 1;
    attribute mti_svvh_generic_type of REG_ADDNSUB1_0_RST : constant is 1;
    attribute mti_svvh_generic_type of REG_ADDNSUB1_1_CLK : constant is 1;
    attribute mti_svvh_generic_type of REG_ADDNSUB1_1_CE : constant is 1;
    attribute mti_svvh_generic_type of REG_ADDNSUB1_1_RST : constant is 1;
    attribute mti_svvh_generic_type of REG_ADDNSUB3_0_CLK : constant is 1;
    attribute mti_svvh_generic_type of REG_ADDNSUB3_0_CE : constant is 1;
    attribute mti_svvh_generic_type of REG_ADDNSUB3_0_RST : constant is 1;
    attribute mti_svvh_generic_type of REG_ADDNSUB3_1_CLK : constant is 1;
    attribute mti_svvh_generic_type of REG_ADDNSUB3_1_CE : constant is 1;
    attribute mti_svvh_generic_type of REG_ADDNSUB3_1_RST : constant is 1;
    attribute mti_svvh_generic_type of GSR : constant is 1;
end MULT18X18ADDSUBSUMB;
