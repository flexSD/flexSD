library verilog;
use verilog.vl_types.all;
entity MULT36X36B is
    generic(
        REG_INPUTA_CLK  : string  := "NONE";
        REG_INPUTA_CE   : string  := "CE0";
        REG_INPUTA_RST  : string  := "RST0";
        REG_INPUTB_CLK  : string  := "NONE";
        REG_INPUTB_CE   : string  := "CE0";
        REG_INPUTB_RST  : string  := "RST0";
        REG_PIPELINE_CLK: string  := "NONE";
        REG_PIPELINE_CE : string  := "CE0";
        REG_PIPELINE_RST: string  := "RST0";
        REG_OUTPUT_CLK  : string  := "NONE";
        REG_OUTPUT_CE   : string  := "CE0";
        REG_OUTPUT_RST  : string  := "RST0";
        REG_SIGNEDA_0_CLK: string  := "NONE";
        REG_SIGNEDA_0_CE: string  := "CE0";
        REG_SIGNEDA_0_RST: string  := "RST0";
        REG_SIGNEDA_1_CLK: string  := "NONE";
        REG_SIGNEDA_1_CE: string  := "CE0";
        REG_SIGNEDA_1_RST: string  := "RST0";
        REG_SIGNEDB_0_CLK: string  := "NONE";
        REG_SIGNEDB_0_CE: string  := "CE0";
        REG_SIGNEDB_0_RST: string  := "RST0";
        REG_SIGNEDB_1_CLK: string  := "NONE";
        REG_SIGNEDB_1_CE: string  := "CE0";
        REG_SIGNEDB_1_RST: string  := "RST0";
        GSR             : string  := "ENABLED"
    );
    port(
        P71             : out    vl_logic;
        P70             : out    vl_logic;
        P69             : out    vl_logic;
        P68             : out    vl_logic;
        P67             : out    vl_logic;
        P66             : out    vl_logic;
        P65             : out    vl_logic;
        P64             : out    vl_logic;
        P63             : out    vl_logic;
        P62             : out    vl_logic;
        P61             : out    vl_logic;
        P60             : out    vl_logic;
        P59             : out    vl_logic;
        P58             : out    vl_logic;
        P57             : out    vl_logic;
        P56             : out    vl_logic;
        P55             : out    vl_logic;
        P54             : out    vl_logic;
        P53             : out    vl_logic;
        P52             : out    vl_logic;
        P51             : out    vl_logic;
        P50             : out    vl_logic;
        P49             : out    vl_logic;
        P48             : out    vl_logic;
        P47             : out    vl_logic;
        P46             : out    vl_logic;
        P45             : out    vl_logic;
        P44             : out    vl_logic;
        P43             : out    vl_logic;
        P42             : out    vl_logic;
        P41             : out    vl_logic;
        P40             : out    vl_logic;
        P39             : out    vl_logic;
        P38             : out    vl_logic;
        P37             : out    vl_logic;
        P36             : out    vl_logic;
        P35             : out    vl_logic;
        P34             : out    vl_logic;
        P33             : out    vl_logic;
        P32             : out    vl_logic;
        P31             : out    vl_logic;
        P30             : out    vl_logic;
        P29             : out    vl_logic;
        P28             : out    vl_logic;
        P27             : out    vl_logic;
        P26             : out    vl_logic;
        P25             : out    vl_logic;
        P24             : out    vl_logic;
        P23             : out    vl_logic;
        P22             : out    vl_logic;
        P21             : out    vl_logic;
        P20             : out    vl_logic;
        P19             : out    vl_logic;
        P18             : out    vl_logic;
        P17             : out    vl_logic;
        P16             : out    vl_logic;
        P15             : out    vl_logic;
        P14             : out    vl_logic;
        P13             : out    vl_logic;
        P12             : out    vl_logic;
        P11             : out    vl_logic;
        P10             : out    vl_logic;
        P9              : out    vl_logic;
        P8              : out    vl_logic;
        P7              : out    vl_logic;
        P6              : out    vl_logic;
        P5              : out    vl_logic;
        P4              : out    vl_logic;
        P3              : out    vl_logic;
        P2              : out    vl_logic;
        P1              : out    vl_logic;
        P0              : out    vl_logic;
        A35             : in     vl_logic;
        A34             : in     vl_logic;
        A33             : in     vl_logic;
        A32             : in     vl_logic;
        A31             : in     vl_logic;
        A30             : in     vl_logic;
        A29             : in     vl_logic;
        A28             : in     vl_logic;
        A27             : in     vl_logic;
        A26             : in     vl_logic;
        A25             : in     vl_logic;
        A24             : in     vl_logic;
        A23             : in     vl_logic;
        A22             : in     vl_logic;
        A21             : in     vl_logic;
        A20             : in     vl_logic;
        A19             : in     vl_logic;
        A18             : in     vl_logic;
        A17             : in     vl_logic;
        A16             : in     vl_logic;
        A15             : in     vl_logic;
        A14             : in     vl_logic;
        A13             : in     vl_logic;
        A12             : in     vl_logic;
        A11             : in     vl_logic;
        A10             : in     vl_logic;
        A9              : in     vl_logic;
        A8              : in     vl_logic;
        A7              : in     vl_logic;
        A6              : in     vl_logic;
        A5              : in     vl_logic;
        A4              : in     vl_logic;
        A3              : in     vl_logic;
        A2              : in     vl_logic;
        A1              : in     vl_logic;
        A0              : in     vl_logic;
        B35             : in     vl_logic;
        B34             : in     vl_logic;
        B33             : in     vl_logic;
        B32             : in     vl_logic;
        B31             : in     vl_logic;
        B30             : in     vl_logic;
        B29             : in     vl_logic;
        B28             : in     vl_logic;
        B27             : in     vl_logic;
        B26             : in     vl_logic;
        B25             : in     vl_logic;
        B24             : in     vl_logic;
        B23             : in     vl_logic;
        B22             : in     vl_logic;
        B21             : in     vl_logic;
        B20             : in     vl_logic;
        B19             : in     vl_logic;
        B18             : in     vl_logic;
        B17             : in     vl_logic;
        B16             : in     vl_logic;
        B15             : in     vl_logic;
        B14             : in     vl_logic;
        B13             : in     vl_logic;
        B12             : in     vl_logic;
        B11             : in     vl_logic;
        B10             : in     vl_logic;
        B9              : in     vl_logic;
        B8              : in     vl_logic;
        B7              : in     vl_logic;
        B6              : in     vl_logic;
        B5              : in     vl_logic;
        B4              : in     vl_logic;
        B3              : in     vl_logic;
        B2              : in     vl_logic;
        B1              : in     vl_logic;
        B0              : in     vl_logic;
        SIGNEDA         : in     vl_logic;
        SIGNEDB         : in     vl_logic;
        CE0             : in     vl_logic;
        CE1             : in     vl_logic;
        CE2             : in     vl_logic;
        CE3             : in     vl_logic;
        CLK0            : in     vl_logic;
        CLK1            : in     vl_logic;
        CLK2            : in     vl_logic;
        CLK3            : in     vl_logic;
        RST0            : in     vl_logic;
        RST1            : in     vl_logic;
        RST2            : in     vl_logic;
        RST3            : in     vl_logic
    );
end MULT36X36B;
