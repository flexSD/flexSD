library verilog;
use verilog.vl_types.all;
entity MULT9X9B is
    generic(
        REG_INPUTA_CLK  : string  := "NONE";
        REG_INPUTA_CE   : string  := "CE0";
        REG_INPUTA_RST  : string  := "RST0";
        REG_INPUTB_CLK  : string  := "NONE";
        REG_INPUTB_CE   : string  := "CE0";
        REG_INPUTB_RST  : string  := "RST0";
        REG_PIPELINE_CLK: string  := "NONE";
        REG_PIPELINE_CE : string  := "CE0";
        REG_PIPELINE_RST: string  := "RST0";
        REG_OUTPUT_CLK  : string  := "NONE";
        REG_OUTPUT_CE   : string  := "CE0";
        REG_OUTPUT_RST  : string  := "RST0";
        REG_SIGNEDA_CLK : string  := "NONE";
        REG_SIGNEDA_CE  : string  := "CE0";
        REG_SIGNEDA_RST : string  := "RST0";
        REG_SIGNEDB_CLK : string  := "NONE";
        REG_SIGNEDB_CE  : string  := "CE0";
        REG_SIGNEDB_RST : string  := "RST0";
        GSR             : string  := "ENABLED"
    );
    port(
        P17             : out    vl_logic;
        P16             : out    vl_logic;
        P15             : out    vl_logic;
        P14             : out    vl_logic;
        P13             : out    vl_logic;
        P12             : out    vl_logic;
        P11             : out    vl_logic;
        P10             : out    vl_logic;
        P9              : out    vl_logic;
        P8              : out    vl_logic;
        P7              : out    vl_logic;
        P6              : out    vl_logic;
        P5              : out    vl_logic;
        P4              : out    vl_logic;
        P3              : out    vl_logic;
        P2              : out    vl_logic;
        P1              : out    vl_logic;
        P0              : out    vl_logic;
        SROA8           : out    vl_logic;
        SROA7           : out    vl_logic;
        SROA6           : out    vl_logic;
        SROA5           : out    vl_logic;
        SROA4           : out    vl_logic;
        SROA3           : out    vl_logic;
        SROA2           : out    vl_logic;
        SROA1           : out    vl_logic;
        SROA0           : out    vl_logic;
        SROB8           : out    vl_logic;
        SROB7           : out    vl_logic;
        SROB6           : out    vl_logic;
        SROB5           : out    vl_logic;
        SROB4           : out    vl_logic;
        SROB3           : out    vl_logic;
        SROB2           : out    vl_logic;
        SROB1           : out    vl_logic;
        SROB0           : out    vl_logic;
        A8              : in     vl_logic;
        A7              : in     vl_logic;
        A6              : in     vl_logic;
        A5              : in     vl_logic;
        A4              : in     vl_logic;
        A3              : in     vl_logic;
        A2              : in     vl_logic;
        A1              : in     vl_logic;
        A0              : in     vl_logic;
        B8              : in     vl_logic;
        B7              : in     vl_logic;
        B6              : in     vl_logic;
        B5              : in     vl_logic;
        B4              : in     vl_logic;
        B3              : in     vl_logic;
        B2              : in     vl_logic;
        B1              : in     vl_logic;
        B0              : in     vl_logic;
        SRIA8           : in     vl_logic;
        SRIA7           : in     vl_logic;
        SRIA6           : in     vl_logic;
        SRIA5           : in     vl_logic;
        SRIA4           : in     vl_logic;
        SRIA3           : in     vl_logic;
        SRIA2           : in     vl_logic;
        SRIA1           : in     vl_logic;
        SRIA0           : in     vl_logic;
        SRIB8           : in     vl_logic;
        SRIB7           : in     vl_logic;
        SRIB6           : in     vl_logic;
        SRIB5           : in     vl_logic;
        SRIB4           : in     vl_logic;
        SRIB3           : in     vl_logic;
        SRIB2           : in     vl_logic;
        SRIB1           : in     vl_logic;
        SRIB0           : in     vl_logic;
        SIGNEDA         : in     vl_logic;
        SIGNEDB         : in     vl_logic;
        CE0             : in     vl_logic;
        CE1             : in     vl_logic;
        CE2             : in     vl_logic;
        CE3             : in     vl_logic;
        CLK0            : in     vl_logic;
        CLK1            : in     vl_logic;
        CLK2            : in     vl_logic;
        CLK3            : in     vl_logic;
        RST0            : in     vl_logic;
        RST1            : in     vl_logic;
        RST2            : in     vl_logic;
        RST3            : in     vl_logic;
        SOURCEA         : in     vl_logic;
        SOURCEB         : in     vl_logic
    );
end MULT9X9B;
