library verilog;
use verilog.vl_types.all;
entity MULT9X9ADDSUBSUMB is
    generic(
        REG_INPUTA0_CLK : string  := "NONE";
        REG_INPUTA0_CE  : string  := "CE0";
        REG_INPUTA0_RST : string  := "RST0";
        REG_INPUTA1_CLK : string  := "NONE";
        REG_INPUTA1_CE  : string  := "CE0";
        REG_INPUTA1_RST : string  := "RST0";
        REG_INPUTA2_CLK : string  := "NONE";
        REG_INPUTA2_CE  : string  := "CE0";
        REG_INPUTA2_RST : string  := "RST0";
        REG_INPUTA3_CLK : string  := "NONE";
        REG_INPUTA3_CE  : string  := "CE0";
        REG_INPUTA3_RST : string  := "RST0";
        REG_INPUTB0_CLK : string  := "NONE";
        REG_INPUTB0_CE  : string  := "CE0";
        REG_INPUTB0_RST : string  := "RST0";
        REG_INPUTB1_CLK : string  := "NONE";
        REG_INPUTB1_CE  : string  := "CE0";
        REG_INPUTB1_RST : string  := "RST0";
        REG_INPUTB2_CLK : string  := "NONE";
        REG_INPUTB2_CE  : string  := "CE0";
        REG_INPUTB2_RST : string  := "RST0";
        REG_INPUTB3_CLK : string  := "NONE";
        REG_INPUTB3_CE  : string  := "CE0";
        REG_INPUTB3_RST : string  := "RST0";
        REG_PIPELINE0_CLK: string  := "NONE";
        REG_PIPELINE0_CE: string  := "CE0";
        REG_PIPELINE0_RST: string  := "RST0";
        REG_PIPELINE1_CLK: string  := "NONE";
        REG_PIPELINE1_CE: string  := "CE0";
        REG_PIPELINE1_RST: string  := "RST0";
        REG_PIPELINE2_CLK: string  := "NONE";
        REG_PIPELINE2_CE: string  := "CE0";
        REG_PIPELINE2_RST: string  := "RST0";
        REG_PIPELINE3_CLK: string  := "NONE";
        REG_PIPELINE3_CE: string  := "CE0";
        REG_PIPELINE3_RST: string  := "RST0";
        REG_OUTPUT_CLK  : string  := "NONE";
        REG_OUTPUT_CE   : string  := "CE0";
        REG_OUTPUT_RST  : string  := "RST0";
        REG_SIGNEDA_0_CLK: string  := "NONE";
        REG_SIGNEDA_0_CE: string  := "CE0";
        REG_SIGNEDA_0_RST: string  := "RST0";
        REG_SIGNEDA_1_CLK: string  := "NONE";
        REG_SIGNEDA_1_CE: string  := "CE0";
        REG_SIGNEDA_1_RST: string  := "RST0";
        REG_SIGNEDB_0_CLK: string  := "NONE";
        REG_SIGNEDB_0_CE: string  := "CE0";
        REG_SIGNEDB_0_RST: string  := "RST0";
        REG_SIGNEDB_1_CLK: string  := "NONE";
        REG_SIGNEDB_1_CE: string  := "CE0";
        REG_SIGNEDB_1_RST: string  := "RST0";
        REG_ADDNSUB1_0_CLK: string  := "NONE";
        REG_ADDNSUB1_0_CE: string  := "CE0";
        REG_ADDNSUB1_0_RST: string  := "RST0";
        REG_ADDNSUB1_1_CLK: string  := "NONE";
        REG_ADDNSUB1_1_CE: string  := "CE0";
        REG_ADDNSUB1_1_RST: string  := "RST0";
        REG_ADDNSUB3_0_CLK: string  := "NONE";
        REG_ADDNSUB3_0_CE: string  := "CE0";
        REG_ADDNSUB3_0_RST: string  := "RST0";
        REG_ADDNSUB3_1_CLK: string  := "NONE";
        REG_ADDNSUB3_1_CE: string  := "CE0";
        REG_ADDNSUB3_1_RST: string  := "RST0";
        GSR             : string  := "ENABLED"
    );
    port(
        SUM19           : out    vl_logic;
        SUM18           : out    vl_logic;
        SUM17           : out    vl_logic;
        SUM16           : out    vl_logic;
        SUM15           : out    vl_logic;
        SUM14           : out    vl_logic;
        SUM13           : out    vl_logic;
        SUM12           : out    vl_logic;
        SUM11           : out    vl_logic;
        SUM10           : out    vl_logic;
        SUM9            : out    vl_logic;
        SUM8            : out    vl_logic;
        SUM7            : out    vl_logic;
        SUM6            : out    vl_logic;
        SUM5            : out    vl_logic;
        SUM4            : out    vl_logic;
        SUM3            : out    vl_logic;
        SUM2            : out    vl_logic;
        SUM1            : out    vl_logic;
        SUM0            : out    vl_logic;
        SROA8           : out    vl_logic;
        SROA7           : out    vl_logic;
        SROA6           : out    vl_logic;
        SROA5           : out    vl_logic;
        SROA4           : out    vl_logic;
        SROA3           : out    vl_logic;
        SROA2           : out    vl_logic;
        SROA1           : out    vl_logic;
        SROA0           : out    vl_logic;
        SROB8           : out    vl_logic;
        SROB7           : out    vl_logic;
        SROB6           : out    vl_logic;
        SROB5           : out    vl_logic;
        SROB4           : out    vl_logic;
        SROB3           : out    vl_logic;
        SROB2           : out    vl_logic;
        SROB1           : out    vl_logic;
        SROB0           : out    vl_logic;
        A08             : in     vl_logic;
        A07             : in     vl_logic;
        A06             : in     vl_logic;
        A05             : in     vl_logic;
        A04             : in     vl_logic;
        A03             : in     vl_logic;
        A02             : in     vl_logic;
        A01             : in     vl_logic;
        A00             : in     vl_logic;
        A18             : in     vl_logic;
        A17             : in     vl_logic;
        A16             : in     vl_logic;
        A15             : in     vl_logic;
        A14             : in     vl_logic;
        A13             : in     vl_logic;
        A12             : in     vl_logic;
        A11             : in     vl_logic;
        A10             : in     vl_logic;
        A28             : in     vl_logic;
        A27             : in     vl_logic;
        A26             : in     vl_logic;
        A25             : in     vl_logic;
        A24             : in     vl_logic;
        A23             : in     vl_logic;
        A22             : in     vl_logic;
        A21             : in     vl_logic;
        A20             : in     vl_logic;
        A38             : in     vl_logic;
        A37             : in     vl_logic;
        A36             : in     vl_logic;
        A35             : in     vl_logic;
        A34             : in     vl_logic;
        A33             : in     vl_logic;
        A32             : in     vl_logic;
        A31             : in     vl_logic;
        A30             : in     vl_logic;
        B08             : in     vl_logic;
        B07             : in     vl_logic;
        B06             : in     vl_logic;
        B05             : in     vl_logic;
        B04             : in     vl_logic;
        B03             : in     vl_logic;
        B02             : in     vl_logic;
        B01             : in     vl_logic;
        B00             : in     vl_logic;
        B18             : in     vl_logic;
        B17             : in     vl_logic;
        B16             : in     vl_logic;
        B15             : in     vl_logic;
        B14             : in     vl_logic;
        B13             : in     vl_logic;
        B12             : in     vl_logic;
        B11             : in     vl_logic;
        B10             : in     vl_logic;
        B28             : in     vl_logic;
        B27             : in     vl_logic;
        B26             : in     vl_logic;
        B25             : in     vl_logic;
        B24             : in     vl_logic;
        B23             : in     vl_logic;
        B22             : in     vl_logic;
        B21             : in     vl_logic;
        B20             : in     vl_logic;
        B38             : in     vl_logic;
        B37             : in     vl_logic;
        B36             : in     vl_logic;
        B35             : in     vl_logic;
        B34             : in     vl_logic;
        B33             : in     vl_logic;
        B32             : in     vl_logic;
        B31             : in     vl_logic;
        B30             : in     vl_logic;
        SRIA8           : in     vl_logic;
        SRIA7           : in     vl_logic;
        SRIA6           : in     vl_logic;
        SRIA5           : in     vl_logic;
        SRIA4           : in     vl_logic;
        SRIA3           : in     vl_logic;
        SRIA2           : in     vl_logic;
        SRIA1           : in     vl_logic;
        SRIA0           : in     vl_logic;
        SRIB8           : in     vl_logic;
        SRIB7           : in     vl_logic;
        SRIB6           : in     vl_logic;
        SRIB5           : in     vl_logic;
        SRIB4           : in     vl_logic;
        SRIB3           : in     vl_logic;
        SRIB2           : in     vl_logic;
        SRIB1           : in     vl_logic;
        SRIB0           : in     vl_logic;
        SIGNEDA         : in     vl_logic;
        SIGNEDB         : in     vl_logic;
        ADDNSUB1        : in     vl_logic;
        ADDNSUB3        : in     vl_logic;
        CE0             : in     vl_logic;
        CE1             : in     vl_logic;
        CE2             : in     vl_logic;
        CE3             : in     vl_logic;
        CLK0            : in     vl_logic;
        CLK1            : in     vl_logic;
        CLK2            : in     vl_logic;
        CLK3            : in     vl_logic;
        RST0            : in     vl_logic;
        RST1            : in     vl_logic;
        RST2            : in     vl_logic;
        RST3            : in     vl_logic;
        SOURCEA0        : in     vl_logic;
        SOURCEA1        : in     vl_logic;
        SOURCEA2        : in     vl_logic;
        SOURCEA3        : in     vl_logic;
        SOURCEB0        : in     vl_logic;
        SOURCEB1        : in     vl_logic;
        SOURCEB2        : in     vl_logic;
        SOURCEB3        : in     vl_logic
    );
end MULT9X9ADDSUBSUMB;
