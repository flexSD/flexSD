library verilog;
use verilog.vl_types.all;
entity VLO is
    port(
        Z               : out    vl_logic
    );
end VLO;
