library verilog;
use verilog.vl_types.all;
entity SDPRAMC is
    generic(
        GSR             : string  := "ENABLED";
        SRMODE          : string  := "LSR_OVER_CE";
        M1MUX           : string  := "VLO";
        M0MUX           : string  := "VLO";
        LSRMUX          : string  := "VLO";
        CEMUX           : string  := "VLO";
        CLKMUX          : string  := "VLO";
        REG1_SD         : string  := "VLO";
        REG0_SD         : string  := "VLO";
        REG1_REGSET     : string  := "RESET";
        REG0_REGSET     : string  := "RESET";
        LSRONMUX        : string  := "LSRMUX";
        initval         : integer := 0;
        XON             : integer := 0;
        CHECK_RAD0      : integer := 0;
        CHECK_RAD1      : integer := 0;
        CHECK_RAD2      : integer := 0;
        CHECK_RAD3      : integer := 0;
        CHECK_WD1       : integer := 0;
        CHECK_WD0       : integer := 0;
        CHECK_WAD0      : integer := 0;
        CHECK_WAD1      : integer := 0;
        CHECK_WAD2      : integer := 0;
        CHECK_WAD3      : integer := 0;
        CHECK_WRE       : integer := 0;
        CHECK_CE        : integer := 0;
        CHECK_LSR       : integer := 0;
        CHECK_M1        : integer := 0;
        CHECK_DI1       : integer := 0;
        CHECK_DI0       : integer := 0;
        CHECK_M0        : integer := 0
    );
    port(
        M1              : in     vl_logic;
        RAD0            : in     vl_logic;
        RAD1            : in     vl_logic;
        RAD2            : in     vl_logic;
        RAD3            : in     vl_logic;
        WD1             : in     vl_logic;
        WD0             : in     vl_logic;
        WAD0            : in     vl_logic;
        WAD1            : in     vl_logic;
        WAD2            : in     vl_logic;
        WAD3            : in     vl_logic;
        WRE             : in     vl_logic;
        WCK             : in     vl_logic;
        M0              : in     vl_logic;
        DI1             : in     vl_logic;
        DI0             : in     vl_logic;
        CE              : in     vl_logic;
        CLK             : in     vl_logic;
        LSR             : in     vl_logic;
        F0              : out    vl_logic;
        Q0              : out    vl_logic;
        F1              : out    vl_logic;
        Q1              : out    vl_logic
    );
end SDPRAMC;
