library verilog;
use verilog.vl_types.all;
entity MULT18X18MACB is
    generic(
        REG_INPUTA_CLK  : string  := "NONE";
        REG_INPUTA_CE   : string  := "CE0";
        REG_INPUTA_RST  : string  := "RST0";
        REG_INPUTB_CLK  : string  := "NONE";
        REG_INPUTB_CE   : string  := "CE0";
        REG_INPUTB_RST  : string  := "RST0";
        REG_PIPELINE_CLK: string  := "NONE";
        REG_PIPELINE_CE : string  := "CE0";
        REG_PIPELINE_RST: string  := "RST0";
        REG_OUTPUT_CLK  : string  := "NONE";
        REG_OUTPUT_CE   : string  := "CE0";
        REG_OUTPUT_RST  : string  := "RST0";
        REG_SIGNEDA_0_CLK: string  := "NONE";
        REG_SIGNEDA_0_CE: string  := "CE0";
        REG_SIGNEDA_0_RST: string  := "RST0";
        REG_SIGNEDA_1_CLK: string  := "NONE";
        REG_SIGNEDA_1_CE: string  := "CE0";
        REG_SIGNEDA_1_RST: string  := "RST0";
        REG_SIGNEDB_0_CLK: string  := "NONE";
        REG_SIGNEDB_0_CE: string  := "CE0";
        REG_SIGNEDB_0_RST: string  := "RST0";
        REG_SIGNEDB_1_CLK: string  := "NONE";
        REG_SIGNEDB_1_CE: string  := "CE0";
        REG_SIGNEDB_1_RST: string  := "RST0";
        REG_ACCUMSLOAD_0_CLK: string  := "NONE";
        REG_ACCUMSLOAD_0_CE: string  := "CE0";
        REG_ACCUMSLOAD_0_RST: string  := "RST0";
        REG_ACCUMSLOAD_1_CLK: string  := "NONE";
        REG_ACCUMSLOAD_1_CE: string  := "CE0";
        REG_ACCUMSLOAD_1_RST: string  := "RST0";
        REG_ADDNSUB_0_CLK: string  := "NONE";
        REG_ADDNSUB_0_CE: string  := "CE0";
        REG_ADDNSUB_0_RST: string  := "RST0";
        REG_ADDNSUB_1_CLK: string  := "NONE";
        REG_ADDNSUB_1_CE: string  := "CE0";
        REG_ADDNSUB_1_RST: string  := "RST0";
        GSR             : string  := "ENABLED"
    );
    port(
        ACCUM51         : out    vl_logic;
        ACCUM50         : out    vl_logic;
        ACCUM49         : out    vl_logic;
        ACCUM48         : out    vl_logic;
        ACCUM47         : out    vl_logic;
        ACCUM46         : out    vl_logic;
        ACCUM45         : out    vl_logic;
        ACCUM44         : out    vl_logic;
        ACCUM43         : out    vl_logic;
        ACCUM42         : out    vl_logic;
        ACCUM41         : out    vl_logic;
        ACCUM40         : out    vl_logic;
        ACCUM39         : out    vl_logic;
        ACCUM38         : out    vl_logic;
        ACCUM37         : out    vl_logic;
        ACCUM36         : out    vl_logic;
        ACCUM35         : out    vl_logic;
        ACCUM34         : out    vl_logic;
        ACCUM33         : out    vl_logic;
        ACCUM32         : out    vl_logic;
        ACCUM31         : out    vl_logic;
        ACCUM30         : out    vl_logic;
        ACCUM29         : out    vl_logic;
        ACCUM28         : out    vl_logic;
        ACCUM27         : out    vl_logic;
        ACCUM26         : out    vl_logic;
        ACCUM25         : out    vl_logic;
        ACCUM24         : out    vl_logic;
        ACCUM23         : out    vl_logic;
        ACCUM22         : out    vl_logic;
        ACCUM21         : out    vl_logic;
        ACCUM20         : out    vl_logic;
        ACCUM19         : out    vl_logic;
        ACCUM18         : out    vl_logic;
        ACCUM17         : out    vl_logic;
        ACCUM16         : out    vl_logic;
        ACCUM15         : out    vl_logic;
        ACCUM14         : out    vl_logic;
        ACCUM13         : out    vl_logic;
        ACCUM12         : out    vl_logic;
        ACCUM11         : out    vl_logic;
        ACCUM10         : out    vl_logic;
        ACCUM9          : out    vl_logic;
        ACCUM8          : out    vl_logic;
        ACCUM7          : out    vl_logic;
        ACCUM6          : out    vl_logic;
        ACCUM5          : out    vl_logic;
        ACCUM4          : out    vl_logic;
        ACCUM3          : out    vl_logic;
        ACCUM2          : out    vl_logic;
        ACCUM1          : out    vl_logic;
        ACCUM0          : out    vl_logic;
        SROA17          : out    vl_logic;
        SROA16          : out    vl_logic;
        SROA15          : out    vl_logic;
        SROA14          : out    vl_logic;
        SROA13          : out    vl_logic;
        SROA12          : out    vl_logic;
        SROA11          : out    vl_logic;
        SROA10          : out    vl_logic;
        SROA9           : out    vl_logic;
        SROA8           : out    vl_logic;
        SROA7           : out    vl_logic;
        SROA6           : out    vl_logic;
        SROA5           : out    vl_logic;
        SROA4           : out    vl_logic;
        SROA3           : out    vl_logic;
        SROA2           : out    vl_logic;
        SROA1           : out    vl_logic;
        SROA0           : out    vl_logic;
        SROB17          : out    vl_logic;
        SROB16          : out    vl_logic;
        SROB15          : out    vl_logic;
        SROB14          : out    vl_logic;
        SROB13          : out    vl_logic;
        SROB12          : out    vl_logic;
        SROB11          : out    vl_logic;
        SROB10          : out    vl_logic;
        SROB9           : out    vl_logic;
        SROB8           : out    vl_logic;
        SROB7           : out    vl_logic;
        SROB6           : out    vl_logic;
        SROB5           : out    vl_logic;
        SROB4           : out    vl_logic;
        SROB3           : out    vl_logic;
        SROB2           : out    vl_logic;
        SROB1           : out    vl_logic;
        SROB0           : out    vl_logic;
        OVERFLOW        : out    vl_logic;
        A17             : in     vl_logic;
        A16             : in     vl_logic;
        A15             : in     vl_logic;
        A14             : in     vl_logic;
        A13             : in     vl_logic;
        A12             : in     vl_logic;
        A11             : in     vl_logic;
        A10             : in     vl_logic;
        A9              : in     vl_logic;
        A8              : in     vl_logic;
        A7              : in     vl_logic;
        A6              : in     vl_logic;
        A5              : in     vl_logic;
        A4              : in     vl_logic;
        A3              : in     vl_logic;
        A2              : in     vl_logic;
        A1              : in     vl_logic;
        A0              : in     vl_logic;
        B17             : in     vl_logic;
        B16             : in     vl_logic;
        B15             : in     vl_logic;
        B14             : in     vl_logic;
        B13             : in     vl_logic;
        B12             : in     vl_logic;
        B11             : in     vl_logic;
        B10             : in     vl_logic;
        B9              : in     vl_logic;
        B8              : in     vl_logic;
        B7              : in     vl_logic;
        B6              : in     vl_logic;
        B5              : in     vl_logic;
        B4              : in     vl_logic;
        B3              : in     vl_logic;
        B2              : in     vl_logic;
        B1              : in     vl_logic;
        B0              : in     vl_logic;
        SRIA17          : in     vl_logic;
        SRIA16          : in     vl_logic;
        SRIA15          : in     vl_logic;
        SRIA14          : in     vl_logic;
        SRIA13          : in     vl_logic;
        SRIA12          : in     vl_logic;
        SRIA11          : in     vl_logic;
        SRIA10          : in     vl_logic;
        SRIA9           : in     vl_logic;
        SRIA8           : in     vl_logic;
        SRIA7           : in     vl_logic;
        SRIA6           : in     vl_logic;
        SRIA5           : in     vl_logic;
        SRIA4           : in     vl_logic;
        SRIA3           : in     vl_logic;
        SRIA2           : in     vl_logic;
        SRIA1           : in     vl_logic;
        SRIA0           : in     vl_logic;
        SRIB17          : in     vl_logic;
        SRIB16          : in     vl_logic;
        SRIB15          : in     vl_logic;
        SRIB14          : in     vl_logic;
        SRIB13          : in     vl_logic;
        SRIB12          : in     vl_logic;
        SRIB11          : in     vl_logic;
        SRIB10          : in     vl_logic;
        SRIB9           : in     vl_logic;
        SRIB8           : in     vl_logic;
        SRIB7           : in     vl_logic;
        SRIB6           : in     vl_logic;
        SRIB5           : in     vl_logic;
        SRIB4           : in     vl_logic;
        SRIB3           : in     vl_logic;
        SRIB2           : in     vl_logic;
        SRIB1           : in     vl_logic;
        SRIB0           : in     vl_logic;
        ADDNSUB         : in     vl_logic;
        SIGNEDA         : in     vl_logic;
        SIGNEDB         : in     vl_logic;
        ACCUMSLOAD      : in     vl_logic;
        CE0             : in     vl_logic;
        CE1             : in     vl_logic;
        CE2             : in     vl_logic;
        CE3             : in     vl_logic;
        CLK0            : in     vl_logic;
        CLK1            : in     vl_logic;
        CLK2            : in     vl_logic;
        CLK3            : in     vl_logic;
        RST0            : in     vl_logic;
        RST1            : in     vl_logic;
        RST2            : in     vl_logic;
        RST3            : in     vl_logic;
        SOURCEA         : in     vl_logic;
        SOURCEB         : in     vl_logic;
        LD51            : in     vl_logic;
        LD50            : in     vl_logic;
        LD49            : in     vl_logic;
        LD48            : in     vl_logic;
        LD47            : in     vl_logic;
        LD46            : in     vl_logic;
        LD45            : in     vl_logic;
        LD44            : in     vl_logic;
        LD43            : in     vl_logic;
        LD42            : in     vl_logic;
        LD41            : in     vl_logic;
        LD40            : in     vl_logic;
        LD39            : in     vl_logic;
        LD38            : in     vl_logic;
        LD37            : in     vl_logic;
        LD36            : in     vl_logic;
        LD35            : in     vl_logic;
        LD34            : in     vl_logic;
        LD33            : in     vl_logic;
        LD32            : in     vl_logic;
        LD31            : in     vl_logic;
        LD30            : in     vl_logic;
        LD29            : in     vl_logic;
        LD28            : in     vl_logic;
        LD27            : in     vl_logic;
        LD26            : in     vl_logic;
        LD25            : in     vl_logic;
        LD24            : in     vl_logic;
        LD23            : in     vl_logic;
        LD22            : in     vl_logic;
        LD21            : in     vl_logic;
        LD20            : in     vl_logic;
        LD19            : in     vl_logic;
        LD18            : in     vl_logic;
        LD17            : in     vl_logic;
        LD16            : in     vl_logic;
        LD15            : in     vl_logic;
        LD14            : in     vl_logic;
        LD13            : in     vl_logic;
        LD12            : in     vl_logic;
        LD11            : in     vl_logic;
        LD10            : in     vl_logic;
        LD9             : in     vl_logic;
        LD8             : in     vl_logic;
        LD7             : in     vl_logic;
        LD6             : in     vl_logic;
        LD5             : in     vl_logic;
        LD4             : in     vl_logic;
        LD3             : in     vl_logic;
        LD2             : in     vl_logic;
        LD1             : in     vl_logic;
        LD0             : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of REG_INPUTA_CLK : constant is 1;
    attribute mti_svvh_generic_type of REG_INPUTA_CE : constant is 1;
    attribute mti_svvh_generic_type of REG_INPUTA_RST : constant is 1;
    attribute mti_svvh_generic_type of REG_INPUTB_CLK : constant is 1;
    attribute mti_svvh_generic_type of REG_INPUTB_CE : constant is 1;
    attribute mti_svvh_generic_type of REG_INPUTB_RST : constant is 1;
    attribute mti_svvh_generic_type of REG_PIPELINE_CLK : constant is 1;
    attribute mti_svvh_generic_type of REG_PIPELINE_CE : constant is 1;
    attribute mti_svvh_generic_type of REG_PIPELINE_RST : constant is 1;
    attribute mti_svvh_generic_type of REG_OUTPUT_CLK : constant is 1;
    attribute mti_svvh_generic_type of REG_OUTPUT_CE : constant is 1;
    attribute mti_svvh_generic_type of REG_OUTPUT_RST : constant is 1;
    attribute mti_svvh_generic_type of REG_SIGNEDA_0_CLK : constant is 1;
    attribute mti_svvh_generic_type of REG_SIGNEDA_0_CE : constant is 1;
    attribute mti_svvh_generic_type of REG_SIGNEDA_0_RST : constant is 1;
    attribute mti_svvh_generic_type of REG_SIGNEDA_1_CLK : constant is 1;
    attribute mti_svvh_generic_type of REG_SIGNEDA_1_CE : constant is 1;
    attribute mti_svvh_generic_type of REG_SIGNEDA_1_RST : constant is 1;
    attribute mti_svvh_generic_type of REG_SIGNEDB_0_CLK : constant is 1;
    attribute mti_svvh_generic_type of REG_SIGNEDB_0_CE : constant is 1;
    attribute mti_svvh_generic_type of REG_SIGNEDB_0_RST : constant is 1;
    attribute mti_svvh_generic_type of REG_SIGNEDB_1_CLK : constant is 1;
    attribute mti_svvh_generic_type of REG_SIGNEDB_1_CE : constant is 1;
    attribute mti_svvh_generic_type of REG_SIGNEDB_1_RST : constant is 1;
    attribute mti_svvh_generic_type of REG_ACCUMSLOAD_0_CLK : constant is 1;
    attribute mti_svvh_generic_type of REG_ACCUMSLOAD_0_CE : constant is 1;
    attribute mti_svvh_generic_type of REG_ACCUMSLOAD_0_RST : constant is 1;
    attribute mti_svvh_generic_type of REG_ACCUMSLOAD_1_CLK : constant is 1;
    attribute mti_svvh_generic_type of REG_ACCUMSLOAD_1_CE : constant is 1;
    attribute mti_svvh_generic_type of REG_ACCUMSLOAD_1_RST : constant is 1;
    attribute mti_svvh_generic_type of REG_ADDNSUB_0_CLK : constant is 1;
    attribute mti_svvh_generic_type of REG_ADDNSUB_0_CE : constant is 1;
    attribute mti_svvh_generic_type of REG_ADDNSUB_0_RST : constant is 1;
    attribute mti_svvh_generic_type of REG_ADDNSUB_1_CLK : constant is 1;
    attribute mti_svvh_generic_type of REG_ADDNSUB_1_CE : constant is 1;
    attribute mti_svvh_generic_type of REG_ADDNSUB_1_RST : constant is 1;
    attribute mti_svvh_generic_type of GSR : constant is 1;
end MULT18X18MACB;
