library verilog;
use verilog.vl_types.all;
entity wb_resync is
    port(
        wb_rst_i        : in     vl_logic;
        wb_clk_i        : in     vl_logic;
        wbs1_cyc_i      : in     vl_logic;
        wbs1_stb_i      : in     vl_logic;
        wbs1_dat_i      : in     vl_logic_vector(31 downto 0);
        wbs1_dat_o      : out    vl_logic_vector(31 downto 0);
        wbs1_ack_o      : out    vl_logic;
        wbs1_we_i       : in     vl_logic;
        wbs1_adr_i      : in     vl_logic_vector(31 downto 0);
        wbs1_sel_i      : in     vl_logic_vector(3 downto 0);
        wbs2_cyc_i      : in     vl_logic;
        wbs2_stb_i      : in     vl_logic;
        wbs2_dat_i      : in     vl_logic_vector(31 downto 0);
        wbs2_dat_o      : out    vl_logic_vector(31 downto 0);
        wbs2_ack_o      : out    vl_logic;
        wbs2_we_i       : in     vl_logic;
        wbs2_adr_i      : in     vl_logic_vector(31 downto 0);
        wbs2_sel_i      : in     vl_logic_vector(3 downto 0);
        wbs3_cyc_i      : in     vl_logic;
        wbs3_stb_i      : in     vl_logic;
        wbs3_dat_i      : in     vl_logic_vector(31 downto 0);
        wbs3_dat_o      : out    vl_logic_vector(31 downto 0);
        wbs3_ack_o      : out    vl_logic;
        wbs3_we_i       : in     vl_logic;
        wbs3_adr_i      : in     vl_logic_vector(31 downto 0);
        wbs3_sel_i      : in     vl_logic_vector(3 downto 0);
        wbs4_cyc_i      : in     vl_logic;
        wbs4_stb_i      : in     vl_logic;
        wbs4_dat_i      : in     vl_logic_vector(31 downto 0);
        wbs4_dat_o      : out    vl_logic_vector(31 downto 0);
        wbs4_ack_o      : out    vl_logic;
        wbs4_we_i       : in     vl_logic;
        wbs4_adr_i      : in     vl_logic_vector(31 downto 0);
        wbs4_sel_i      : in     vl_logic_vector(3 downto 0);
        wbm_clk_i       : in     vl_logic;
        wbm_cyc_o       : out    vl_logic;
        wbm_stb_o       : out    vl_logic;
        wbm_adr_o       : out    vl_logic_vector(31 downto 0);
        wbm_dat_o       : out    vl_logic_vector(31 downto 0);
        wbm_ack_i       : in     vl_logic;
        wbm_dat_i       : in     vl_logic_vector(31 downto 0);
        wbm_we_o        : out    vl_logic;
        wbm_sel_o       : out    vl_logic_vector(3 downto 0)
    );
end wb_resync;
