library verilog;
use verilog.vl_types.all;
entity START is
    port(
        STARTCLK        : in     vl_logic
    );
end START;
