library verilog;
use verilog.vl_types.all;
entity SGSR is
    port(
        GSR             : in     vl_logic;
        CLK             : in     vl_logic
    );
end SGSR;
