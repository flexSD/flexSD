library verilog;
use verilog.vl_types.all;
entity IOWAKEUPA is
    port(
        UWKUP           : in     vl_logic
    );
end IOWAKEUPA;
