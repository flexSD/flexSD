library verilog;
use verilog.vl_types.all;
entity IB is
    port(
        I               : in     vl_logic;
        O               : out    vl_logic
    );
end IB;
