module wb_biquad_interface(

	wb_clk_i,
	wb_rst_i,
	
	log_wbm_cyc_o,
	log_wbm_stb_o,
	log_wbm_we_o,
	log_wbm_adr_o,
	log_wbm_dat_o,
	log_wbm_ack_i,
	
	coeff_wbm_cyc_o,
	coeff_wbm_stb_o,
	coeff_wbm_adr_o,
	coeff_wbm_dat_i,
	coeff_wbm_ack_i,
	
	load_new_coefficients,
	done_loading,
	
	sigmaDeltaInput,
	sigmaDeltaOutput,
	
	filter_clk_i

);

//Clock and reset
input wb_clk_i;
input wb_rst_i;

input filter_clk_i;

//Logging BRAM wishbone interface (write only)
output 			log_wbm_cyc_o;
output 			log_wbm_stb_o;
output			log_wbm_we_o;
output 	[11:0]	log_wbm_adr_o;
output	[15:0]	log_wbm_dat_o;
input			log_wbm_ack_i;
	
//Coefficient BRAM wishbone interface (read only)
output			coeff_wbm_cyc_o;
output			coeff_wbm_stb_o;
output	[8:0]	coeff_wbm_adr_o;
input	[63:0]	coeff_wbm_dat_i;
input			coeff_wbm_ack_i;

//Coefficient update signal, done updating signal
input			load_new_coefficients;
output			done_loading;

//Sigma delta streams for input and output of filter(s)
input			sigmaDeltaInput;
output			sigmaDeltaOutput;

//Store initial values for delay blocks in filter
reg 	[31:0]	delay1_ivalue, delay2_ivalue, delay3_ivalue, delay4_ivalue, sdDelay_ivalue;

//State machine variable
reg		[2:0]	load_state;

//Reset signal generated by state machine for biquad
reg				filter_reset;

//Output to tell coefficient memorywindow that coefficient load has completed
reg         	load_done;

//Coefficient storage registers - passed on to biquad filter module
reg		[31:0]	ffGain1, ffGain2, ffGain3, ffGain4, ffGain5;
reg		[31:0]	fbGain1, fbGain2, fbGain3, fbGain4;
//reg		[2:0]	inlineGain1, inlineGain2, inlineGain3, inlineGain4;

//Wishbone connections for coefficient bram communication
reg				coeff_wbm_cyc, coeff_wbm_stb;
reg		[8:0]	coeff_wbm_adr;

//Main state machine to load coefficients into biquad
always@(posedge wb_clk_i) begin
	
	//If wishbone bus resets, all delay values in filter set to zero, and set state variable to zero
	if(wb_rst_i) begin
		
		//Initial delay register values in biquad
		delay1_ivalue <= 0;
		delay2_ivalue <= 0;
		delay3_ivalue <= 0;
		delay4_ivalue <= 0;
		sdDelay_ivalue <= 0;
		
		//Initial coefficient values
		ffGain1 <= 0;
		ffGain2 <= 0;
		ffGain3 <= 0;
		ffGain4 <= 0;
		ffGain5 <= 0;
	
		fbGain1 <= 0;
		fbGain2 <= 0;
		fbGain3 <= 0;
		fbGain4 <= 0;
	
		//inlineGain1 <= 0;
		//inlineGain2 <= 0;
		//inlineGain3 <= 0;
		//inlineGain4 <= 0;
		
		//Initial internal register values
		load_state <= 3'd0;
		load_done <= 1'b1;
		filter_reset <= 1'b0;
		
	end
	
	//Coefficient load state machine
	case(load_state)
		
		3'd0: begin				
					
			//Run through state machine again when load coefficient wire is asserted
			if(load_new_coefficients) begin
				load_state <= 3'd1;
				load_done <= 1'b0;				//Assert load in progress
			end
		end
			
		3'd1: begin				
			//Begin wb cycle, address 1st 64 bits of coefficient bram
			coeff_wbm_cyc <= 1'b1;
			coeff_wbm_stb <= 1'b1;
			coeff_wbm_adr <= 9'd0;
		
			//When ack is rx'ed, load data from bus into coefficient register and end bus cycle, move to next state
			if(coeff_wbm_ack_i) begin					
				ffGain1 <= coeff_wbm_dat_i[31:0];
				ffGain2 <= coeff_wbm_dat_i[63:32];
				
				coeff_wbm_cyc <= 1'b0;
				coeff_wbm_stb <= 1'b0;
				
				load_state <= 3'd2;	
			end				
		end
		
		3'd2: begin				
			//Begin wb cycle, address 2nd 64 bits of coefficient bram
			coeff_wbm_cyc <= 1'b1;
			coeff_wbm_stb <= 1'b1;
			coeff_wbm_adr <= 9'd1;
			
			//When ack is rx'ed, load data from bus into coefficient register and end bus cycle, move to next state
			if(coeff_wbm_ack_i) begin					
				ffGain3 <= coeff_wbm_dat_i[31:0];
				ffGain4 <= coeff_wbm_dat_i[63:32];
				
				coeff_wbm_cyc <= 1'b0;
				coeff_wbm_stb <= 1'b0;
				
				load_state <= 3'd3;					
			end				
		end
		
		3'd3: begin				
			//Begin wb cycle, address 3rd 64 bits of coefficient bram
			coeff_wbm_cyc <= 1'b1;
			coeff_wbm_stb <= 1'b1;
			coeff_wbm_adr <= 9'd2;
			
			//When ack is rx'ed, load data from bus into coefficient register and end bus cycle, move to next state
			if(coeff_wbm_ack_i) begin					
				ffGain5 <= coeff_wbm_dat_i[31:0];
				fbGain1 <= coeff_wbm_dat_i[63:32];
				
				coeff_wbm_cyc <= 1'b0;
				coeff_wbm_stb <= 1'b0;
				
				load_state <= 3'd4;	
			end				
		end
		
		3'd4: begin				
			//Begin wb cycle, address 4th 64 bits of coefficient bram
			coeff_wbm_cyc <= 1'b1;
			coeff_wbm_stb <= 1'b1;
			coeff_wbm_adr <= 9'd3;
			
			//When ack is rx'ed, load data from bus into coefficient register and end bus cycle, move to next state
			if(coeff_wbm_ack_i) begin					
				fbGain2 <= coeff_wbm_dat_i[31:0];
				fbGain3 <= coeff_wbm_dat_i[63:32];
				
				coeff_wbm_cyc <= 1'b0;
				coeff_wbm_stb <= 1'b0;
				
				load_state <= 3'd5;	
			end				
		end
		
		3'd5: begin				
			//Begin wb cycle, address 5th 64 bits of coefficient bram
			coeff_wbm_cyc <= 1'b1;
			coeff_wbm_stb <= 1'b1;
			coeff_wbm_adr <= 9'd4;
			
			//When ack is rx'ed, load data from bus into coefficient register and end bus cycle, move to idle state
			if(coeff_wbm_ack_i) begin					
				fbGain4 <= coeff_wbm_dat_i[31:0];
				
				//inlineGain1 <= coeff_wbm_dat_i[34:32];
				//inlineGain2 <= coeff_wbm_dat_i[37:35];
				//inlineGain3 <= coeff_wbm_dat_i[40:38];
				//inlineGain4 <= coeff_wbm_dat_i[43:41];
				
				coeff_wbm_cyc <= 1'b0;
				coeff_wbm_stb <= 1'b0;
				
				load_done <= 1'b1;		//Assert to memory window that the coefficient load is done
				
				filter_reset <= 1'b1;		//Reset biquad, loads initial values into delay blocks (required to preserve previous filter state when time multiplexing)
								
				load_state <= 3'd6;
			end				
		end
		
		3'd6: begin
			filter_reset <= 1'b0;			//Reset high for one clock cycle
			load_state <= 3'd0;				//Back to idle state
		end
	
	endcase
	
end

assign coeff_wbm_cyc_o = coeff_wbm_cyc;
assign coeff_wbm_stb_o = coeff_wbm_stb;
assign coeff_wbm_adr_o = coeff_wbm_adr;
assign done_loading = load_done;

biquad_filter_32bit #(0) biquad(	//Loading constant bit shift as parameter

	.filter_clock(filter_clk_i),// && filter_clock_en),
	.reset(filter_reset),

	.mainIn(sigmaDeltaInput),
	.mainOut(sigmaDeltaOutput),
	
	.ffGain1(ffGain1),
	.ffGain2(ffGain2),
	.ffGain3(ffGain3),
	.ffGain4(ffGain4),
	.ffGain5(ffGain5),
	
	.fbGain1(fbGain1),
	.fbGain2(fbGain2),
	.fbGain3(fbGain3),
	.fbGain4(fbGain4),
	
	//.inlineGain1(inlineGain1),
	//.inlineGain2(inlineGain2),
	//.inlineGain3(inlineGain3),
	//.inlineGain4(inlineGain4),
	
	.delay1_ivalue(delay1_ivalue),
	.delay2_ivalue(delay2_ivalue),
	.delay3_ivalue(delay3_ivalue),
	.delay4_ivalue(delay4_ivalue),
	.sdDelay_ivalue(sdDelay_ivalue)

);

endmodule