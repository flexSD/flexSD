library verilog;
use verilog.vl_types.all;
entity slice_tb is
    generic(
        input_bitwidth  : integer := 24
    );
end slice_tb;
