module peripheral_control(

	clk25,
	wb_rst,

	// Hardware Pins
	spi_dat,
	dac_cs,
	
	pga_dat,
	pga_clk,
	
	shiftreg_clr,
	shiftreg_outputreg_clk

);