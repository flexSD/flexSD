library verilog;
use verilog.vl_types.all;
entity PDPW16KB is
    generic(
        DATA_WIDTH_W    : integer := 36;
        DATA_WIDTH_R    : integer := 36;
        REGMODE         : string  := "NOREG";
        RESETMODE       : string  := "SYNC";
        CSDECODE_W      : integer := 0;
        CSDECODE_R      : integer := 0;
        GSR             : string  := "DISABLED";
        INITVAL_00      : integer := 0;
        INITVAL_01      : integer := 0;
        INITVAL_02      : integer := 0;
        INITVAL_03      : integer := 0;
        INITVAL_04      : integer := 0;
        INITVAL_05      : integer := 0;
        INITVAL_06      : integer := 0;
        INITVAL_07      : integer := 0;
        INITVAL_08      : integer := 0;
        INITVAL_09      : integer := 0;
        INITVAL_0A      : integer := 0;
        INITVAL_0B      : integer := 0;
        INITVAL_0C      : integer := 0;
        INITVAL_0D      : integer := 0;
        INITVAL_0E      : integer := 0;
        INITVAL_0F      : integer := 0;
        INITVAL_10      : integer := 0;
        INITVAL_11      : integer := 0;
        INITVAL_12      : integer := 0;
        INITVAL_13      : integer := 0;
        INITVAL_14      : integer := 0;
        INITVAL_15      : integer := 0;
        INITVAL_16      : integer := 0;
        INITVAL_17      : integer := 0;
        INITVAL_18      : integer := 0;
        INITVAL_19      : integer := 0;
        INITVAL_1A      : integer := 0;
        INITVAL_1B      : integer := 0;
        INITVAL_1C      : integer := 0;
        INITVAL_1D      : integer := 0;
        INITVAL_1E      : integer := 0;
        INITVAL_1F      : integer := 0;
        INITVAL_20      : integer := 0;
        INITVAL_21      : integer := 0;
        INITVAL_22      : integer := 0;
        INITVAL_23      : integer := 0;
        INITVAL_24      : integer := 0;
        INITVAL_25      : integer := 0;
        INITVAL_26      : integer := 0;
        INITVAL_27      : integer := 0;
        INITVAL_28      : integer := 0;
        INITVAL_29      : integer := 0;
        INITVAL_2A      : integer := 0;
        INITVAL_2B      : integer := 0;
        INITVAL_2C      : integer := 0;
        INITVAL_2D      : integer := 0;
        INITVAL_2E      : integer := 0;
        INITVAL_2F      : integer := 0;
        INITVAL_30      : integer := 0;
        INITVAL_31      : integer := 0;
        INITVAL_32      : integer := 0;
        INITVAL_33      : integer := 0;
        INITVAL_34      : integer := 0;
        INITVAL_35      : integer := 0;
        INITVAL_36      : integer := 0;
        INITVAL_37      : integer := 0;
        INITVAL_38      : integer := 0;
        INITVAL_39      : integer := 0;
        INITVAL_3A      : integer := 0;
        INITVAL_3B      : integer := 0;
        INITVAL_3C      : integer := 0;
        INITVAL_3D      : integer := 0;
        INITVAL_3E      : integer := 0;
        INITVAL_3F      : integer := 0
    );
    port(
        DI0             : in     vl_logic;
        DI1             : in     vl_logic;
        DI2             : in     vl_logic;
        DI3             : in     vl_logic;
        DI4             : in     vl_logic;
        DI5             : in     vl_logic;
        DI6             : in     vl_logic;
        DI7             : in     vl_logic;
        DI8             : in     vl_logic;
        DI9             : in     vl_logic;
        DI10            : in     vl_logic;
        DI11            : in     vl_logic;
        DI12            : in     vl_logic;
        DI13            : in     vl_logic;
        DI14            : in     vl_logic;
        DI15            : in     vl_logic;
        DI16            : in     vl_logic;
        DI17            : in     vl_logic;
        DI18            : in     vl_logic;
        DI19            : in     vl_logic;
        DI20            : in     vl_logic;
        DI21            : in     vl_logic;
        DI22            : in     vl_logic;
        DI23            : in     vl_logic;
        DI24            : in     vl_logic;
        DI25            : in     vl_logic;
        DI26            : in     vl_logic;
        DI27            : in     vl_logic;
        DI28            : in     vl_logic;
        DI29            : in     vl_logic;
        DI30            : in     vl_logic;
        DI31            : in     vl_logic;
        DI32            : in     vl_logic;
        DI33            : in     vl_logic;
        DI34            : in     vl_logic;
        DI35            : in     vl_logic;
        ADW0            : in     vl_logic;
        ADW1            : in     vl_logic;
        ADW2            : in     vl_logic;
        ADW3            : in     vl_logic;
        ADW4            : in     vl_logic;
        ADW5            : in     vl_logic;
        ADW6            : in     vl_logic;
        ADW7            : in     vl_logic;
        ADW8            : in     vl_logic;
        BE0             : in     vl_logic;
        BE1             : in     vl_logic;
        BE2             : in     vl_logic;
        BE3             : in     vl_logic;
        CEW             : in     vl_logic;
        CLKW            : in     vl_logic;
        CSW0            : in     vl_logic;
        CSW1            : in     vl_logic;
        CSW2            : in     vl_logic;
        ADR0            : in     vl_logic;
        ADR1            : in     vl_logic;
        ADR2            : in     vl_logic;
        ADR3            : in     vl_logic;
        ADR4            : in     vl_logic;
        ADR5            : in     vl_logic;
        ADR6            : in     vl_logic;
        ADR7            : in     vl_logic;
        ADR8            : in     vl_logic;
        ADR9            : in     vl_logic;
        ADR10           : in     vl_logic;
        ADR11           : in     vl_logic;
        ADR12           : in     vl_logic;
        ADR13           : in     vl_logic;
        CER             : in     vl_logic;
        CLKR            : in     vl_logic;
        CSR0            : in     vl_logic;
        CSR1            : in     vl_logic;
        CSR2            : in     vl_logic;
        RST             : in     vl_logic;
        DO0             : out    vl_logic;
        DO1             : out    vl_logic;
        DO2             : out    vl_logic;
        DO3             : out    vl_logic;
        DO4             : out    vl_logic;
        DO5             : out    vl_logic;
        DO6             : out    vl_logic;
        DO7             : out    vl_logic;
        DO8             : out    vl_logic;
        DO9             : out    vl_logic;
        DO10            : out    vl_logic;
        DO11            : out    vl_logic;
        DO12            : out    vl_logic;
        DO13            : out    vl_logic;
        DO14            : out    vl_logic;
        DO15            : out    vl_logic;
        DO16            : out    vl_logic;
        DO17            : out    vl_logic;
        DO18            : out    vl_logic;
        DO19            : out    vl_logic;
        DO20            : out    vl_logic;
        DO21            : out    vl_logic;
        DO22            : out    vl_logic;
        DO23            : out    vl_logic;
        DO24            : out    vl_logic;
        DO25            : out    vl_logic;
        DO26            : out    vl_logic;
        DO27            : out    vl_logic;
        DO28            : out    vl_logic;
        DO29            : out    vl_logic;
        DO30            : out    vl_logic;
        DO31            : out    vl_logic;
        DO32            : out    vl_logic;
        DO33            : out    vl_logic;
        DO34            : out    vl_logic;
        DO35            : out    vl_logic
    );
end PDPW16KB;
