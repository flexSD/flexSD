library verilog;
use verilog.vl_types.all;
entity VHI is
    port(
        Z               : out    vl_logic
    );
end VHI;
