library verilog;
use verilog.vl_types.all;
entity OBZ is
    port(
        I               : in     vl_logic;
        T               : in     vl_logic;
        O               : out    vl_logic
    );
end OBZ;
