library verilog;
use verilog.vl_types.all;
entity DP16KB is
    generic(
        DATA_WIDTH_A    : integer := 18;
        DATA_WIDTH_B    : integer := 18;
        REGMODE_A       : string  := "NOREG";
        REGMODE_B       : string  := "NOREG";
        RESETMODE       : string  := "SYNC";
        CSDECODE_A      : integer := 0;
        CSDECODE_B      : integer := 0;
        WRITEMODE_A     : string  := "NORMAL";
        WRITEMODE_B     : string  := "NORMAL";
        GSR             : string  := "DISABLED";
        INITVAL_00      : integer := 0;
        INITVAL_01      : integer := 0;
        INITVAL_02      : integer := 0;
        INITVAL_03      : integer := 0;
        INITVAL_04      : integer := 0;
        INITVAL_05      : integer := 0;
        INITVAL_06      : integer := 0;
        INITVAL_07      : integer := 0;
        INITVAL_08      : integer := 0;
        INITVAL_09      : integer := 0;
        INITVAL_0A      : integer := 0;
        INITVAL_0B      : integer := 0;
        INITVAL_0C      : integer := 0;
        INITVAL_0D      : integer := 0;
        INITVAL_0E      : integer := 0;
        INITVAL_0F      : integer := 0;
        INITVAL_10      : integer := 0;
        INITVAL_11      : integer := 0;
        INITVAL_12      : integer := 0;
        INITVAL_13      : integer := 0;
        INITVAL_14      : integer := 0;
        INITVAL_15      : integer := 0;
        INITVAL_16      : integer := 0;
        INITVAL_17      : integer := 0;
        INITVAL_18      : integer := 0;
        INITVAL_19      : integer := 0;
        INITVAL_1A      : integer := 0;
        INITVAL_1B      : integer := 0;
        INITVAL_1C      : integer := 0;
        INITVAL_1D      : integer := 0;
        INITVAL_1E      : integer := 0;
        INITVAL_1F      : integer := 0;
        INITVAL_20      : integer := 0;
        INITVAL_21      : integer := 0;
        INITVAL_22      : integer := 0;
        INITVAL_23      : integer := 0;
        INITVAL_24      : integer := 0;
        INITVAL_25      : integer := 0;
        INITVAL_26      : integer := 0;
        INITVAL_27      : integer := 0;
        INITVAL_28      : integer := 0;
        INITVAL_29      : integer := 0;
        INITVAL_2A      : integer := 0;
        INITVAL_2B      : integer := 0;
        INITVAL_2C      : integer := 0;
        INITVAL_2D      : integer := 0;
        INITVAL_2E      : integer := 0;
        INITVAL_2F      : integer := 0;
        INITVAL_30      : integer := 0;
        INITVAL_31      : integer := 0;
        INITVAL_32      : integer := 0;
        INITVAL_33      : integer := 0;
        INITVAL_34      : integer := 0;
        INITVAL_35      : integer := 0;
        INITVAL_36      : integer := 0;
        INITVAL_37      : integer := 0;
        INITVAL_38      : integer := 0;
        INITVAL_39      : integer := 0;
        INITVAL_3A      : integer := 0;
        INITVAL_3B      : integer := 0;
        INITVAL_3C      : integer := 0;
        INITVAL_3D      : integer := 0;
        INITVAL_3E      : integer := 0;
        INITVAL_3F      : integer := 0
    );
    port(
        DIA0            : in     vl_logic;
        DIA1            : in     vl_logic;
        DIA2            : in     vl_logic;
        DIA3            : in     vl_logic;
        DIA4            : in     vl_logic;
        DIA5            : in     vl_logic;
        DIA6            : in     vl_logic;
        DIA7            : in     vl_logic;
        DIA8            : in     vl_logic;
        DIA9            : in     vl_logic;
        DIA10           : in     vl_logic;
        DIA11           : in     vl_logic;
        DIA12           : in     vl_logic;
        DIA13           : in     vl_logic;
        DIA14           : in     vl_logic;
        DIA15           : in     vl_logic;
        DIA16           : in     vl_logic;
        DIA17           : in     vl_logic;
        ADA0            : in     vl_logic;
        ADA1            : in     vl_logic;
        ADA2            : in     vl_logic;
        ADA3            : in     vl_logic;
        ADA4            : in     vl_logic;
        ADA5            : in     vl_logic;
        ADA6            : in     vl_logic;
        ADA7            : in     vl_logic;
        ADA8            : in     vl_logic;
        ADA9            : in     vl_logic;
        ADA10           : in     vl_logic;
        ADA11           : in     vl_logic;
        ADA12           : in     vl_logic;
        ADA13           : in     vl_logic;
        CEA             : in     vl_logic;
        CLKA            : in     vl_logic;
        WEA             : in     vl_logic;
        CSA0            : in     vl_logic;
        CSA1            : in     vl_logic;
        CSA2            : in     vl_logic;
        RSTA            : in     vl_logic;
        DIB0            : in     vl_logic;
        DIB1            : in     vl_logic;
        DIB2            : in     vl_logic;
        DIB3            : in     vl_logic;
        DIB4            : in     vl_logic;
        DIB5            : in     vl_logic;
        DIB6            : in     vl_logic;
        DIB7            : in     vl_logic;
        DIB8            : in     vl_logic;
        DIB9            : in     vl_logic;
        DIB10           : in     vl_logic;
        DIB11           : in     vl_logic;
        DIB12           : in     vl_logic;
        DIB13           : in     vl_logic;
        DIB14           : in     vl_logic;
        DIB15           : in     vl_logic;
        DIB16           : in     vl_logic;
        DIB17           : in     vl_logic;
        ADB0            : in     vl_logic;
        ADB1            : in     vl_logic;
        ADB2            : in     vl_logic;
        ADB3            : in     vl_logic;
        ADB4            : in     vl_logic;
        ADB5            : in     vl_logic;
        ADB6            : in     vl_logic;
        ADB7            : in     vl_logic;
        ADB8            : in     vl_logic;
        ADB9            : in     vl_logic;
        ADB10           : in     vl_logic;
        ADB11           : in     vl_logic;
        ADB12           : in     vl_logic;
        ADB13           : in     vl_logic;
        CEB             : in     vl_logic;
        CLKB            : in     vl_logic;
        WEB             : in     vl_logic;
        CSB0            : in     vl_logic;
        CSB1            : in     vl_logic;
        CSB2            : in     vl_logic;
        RSTB            : in     vl_logic;
        DOA0            : out    vl_logic;
        DOA1            : out    vl_logic;
        DOA2            : out    vl_logic;
        DOA3            : out    vl_logic;
        DOA4            : out    vl_logic;
        DOA5            : out    vl_logic;
        DOA6            : out    vl_logic;
        DOA7            : out    vl_logic;
        DOA8            : out    vl_logic;
        DOA9            : out    vl_logic;
        DOA10           : out    vl_logic;
        DOA11           : out    vl_logic;
        DOA12           : out    vl_logic;
        DOA13           : out    vl_logic;
        DOA14           : out    vl_logic;
        DOA15           : out    vl_logic;
        DOA16           : out    vl_logic;
        DOA17           : out    vl_logic;
        DOB0            : out    vl_logic;
        DOB1            : out    vl_logic;
        DOB2            : out    vl_logic;
        DOB3            : out    vl_logic;
        DOB4            : out    vl_logic;
        DOB5            : out    vl_logic;
        DOB6            : out    vl_logic;
        DOB7            : out    vl_logic;
        DOB8            : out    vl_logic;
        DOB9            : out    vl_logic;
        DOB10           : out    vl_logic;
        DOB11           : out    vl_logic;
        DOB12           : out    vl_logic;
        DOB13           : out    vl_logic;
        DOB14           : out    vl_logic;
        DOB15           : out    vl_logic;
        DOB16           : out    vl_logic;
        DOB17           : out    vl_logic
    );
end DP16KB;
