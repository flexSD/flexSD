library verilog;
use verilog.vl_types.all;
entity IFS1S1B is
    generic(
        GSR             : string  := "ENABLED"
    );
    port(
        D               : in     vl_logic;
        SCLK            : in     vl_logic;
        PD              : in     vl_logic;
        Q               : out    vl_logic
    );
end IFS1S1B;
