library verilog;
use verilog.vl_types.all;
entity slice_vliw_tb is
    generic(
        input_bitwidth  : integer := 24
    );
end slice_vliw_tb;
