library verilog;
use verilog.vl_types.all;
entity UDFDL1_UDP_X is
    // This module cannot be connected to from
    // VHDL because it has unnamed ports.
end UDFDL1_UDP_X;
