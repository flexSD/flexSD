library verilog;
use verilog.vl_types.all;
entity adder_tb is
    generic(
        input_bitwidth  : integer := 24
    );
end adder_tb;
