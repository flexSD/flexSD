library verilog;
use verilog.vl_types.all;
entity ts7500_top is
    port(
        cpu_clkout_pad  : in     vl_logic;
        fpga_25mhz_pad  : in     vl_logic;
        clk_32khz_pad   : out    vl_logic;
        dio_pad         : inout  vl_logic_vector(40 downto 0);
        cpu_uart_txd_pad: in     vl_logic;
        cpu_uart_rxd_pad: out    vl_logic;
        spi_clk_pad     : in     vl_logic;
        spi_mosi_pad    : in     vl_logic;
        spi_miso_pad    : inout  vl_logic;
        gpio_a0_pad     : out    vl_logic;
        gpio_a1_pad     : out    vl_logic;
        gpio_a13_pad    : inout  vl_logic;
        gpio_a14_pad    : inout  vl_logic;
        gpio_a3_pad     : inout  vl_logic;
        gpio_a15_pad    : inout  vl_logic;
        gpio_a16_pad    : inout  vl_logic;
        gpio_a17_pad    : inout  vl_logic;
        gpio_a28_pad    : inout  vl_logic;
        gpio_a29_pad    : inout  vl_logic;
        int28_pad       : inout  vl_logic;
        gpio_a22_pad    : inout  vl_logic;
        gpio_a23_pad    : inout  vl_logic;
        un_reset_pad    : out    vl_logic;
        wd_resetn_pad   : inout  vl_logic;
        en_sd_power_pad : out    vl_logic;
        sd_d0_pad       : inout  vl_logic;
        sd_d1_pad       : inout  vl_logic;
        sd_d2_pad       : inout  vl_logic;
        sd_d3_pad       : inout  vl_logic;
        sd_cmd_pad      : inout  vl_logic;
        sd_clk_pad      : out    vl_logic;
        red_led_pad     : out    vl_logic;
        green_led_pad   : out    vl_logic;
        eth_left_ledn_pad: out    vl_logic;
        eth_right_ledn_pad: out    vl_logic;
        rtc_sda_pad     : inout  vl_logic;
        rtc_scl_pad     : out    vl_logic;
        rtc_int1_pad    : in     vl_logic;
        ser_flash_wp_padn: out    vl_logic;
        ser_flash_cs_padn: out    vl_logic;
        flash_clk_pad   : out    vl_logic;
        flash_mosi_pad  : out    vl_logic;
        flash_miso_pad  : in     vl_logic
    );
end ts7500_top;
